`timescale 1ns / 1ps
module cos_rom (
    input  logic        [8:0] addr,
    output logic signed [8:0] re,  // 실수부
    output logic signed [8:0] im   // 허수부
);

    // ROM 선언
    wire signed [8:0] rom_re[511:0];
    wire signed [8:0] rom_im[511:0];

    assign re = rom_re[addr];
    assign im = rom_im[addr];

    // cos_rom_re_assign.txt
    assign rom_im[0] = 9'sd0;
    assign rom_im[1] = 9'sd0;
    assign rom_im[2] = 9'sd0;
    assign rom_im[3] = 9'sd0;
    assign rom_im[4] = 9'sd0;
    assign rom_im[5] = 9'sd0;
    assign rom_im[6] = 9'sd0;
    assign rom_im[7] = 9'sd0;
    assign rom_im[8] = 9'sd0;
    assign rom_im[9] = 9'sd0;
    assign rom_im[10] = 9'sd0;
    assign rom_im[11] = 9'sd0;
    assign rom_im[12] = 9'sd0;
    assign rom_im[13] = 9'sd0;
    assign rom_im[14] = 9'sd0;
    assign rom_im[15] = 9'sd0;
    assign rom_im[16] = 9'sd0;
    assign rom_im[17] = 9'sd0;
    assign rom_im[18] = 9'sd0;
    assign rom_im[19] = 9'sd0;
    assign rom_im[20] = 9'sd0;
    assign rom_im[21] = 9'sd0;
    assign rom_im[22] = 9'sd0;
    assign rom_im[23] = 9'sd0;
    assign rom_im[24] = 9'sd0;
    assign rom_im[25] = 9'sd0;
    assign rom_im[26] = 9'sd0;
    assign rom_im[27] = 9'sd0;
    assign rom_im[28] = 9'sd0;
    assign rom_im[29] = 9'sd0;
    assign rom_im[30] = 9'sd0;
    assign rom_im[31] = 9'sd0;
    assign rom_im[32] = 9'sd0;
    assign rom_im[33] = 9'sd0;
    assign rom_im[34] = 9'sd0;
    assign rom_im[35] = 9'sd0;
    assign rom_im[36] = 9'sd0;
    assign rom_im[37] = 9'sd0;
    assign rom_im[38] = 9'sd0;
    assign rom_im[39] = 9'sd0;
    assign rom_im[40] = 9'sd0;
    assign rom_im[41] = 9'sd0;
    assign rom_im[42] = 9'sd0;
    assign rom_im[43] = 9'sd0;
    assign rom_im[44] = 9'sd0;
    assign rom_im[45] = 9'sd0;
    assign rom_im[46] = 9'sd0;
    assign rom_im[47] = 9'sd0;
    assign rom_im[48] = 9'sd0;
    assign rom_im[49] = 9'sd0;
    assign rom_im[50] = 9'sd0;
    assign rom_im[51] = 9'sd0;
    assign rom_im[52] = 9'sd0;
    assign rom_im[53] = 9'sd0;
    assign rom_im[54] = 9'sd0;
    assign rom_im[55] = 9'sd0;
    assign rom_im[56] = 9'sd0;
    assign rom_im[57] = 9'sd0;
    assign rom_im[58] = 9'sd0;
    assign rom_im[59] = 9'sd0;
    assign rom_im[60] = 9'sd0;
    assign rom_im[61] = 9'sd0;
    assign rom_im[62] = 9'sd0;
    assign rom_im[63] = 9'sd0;
    assign rom_im[64] = 9'sd0;
    assign rom_im[65] = 9'sd0;
    assign rom_im[66] = 9'sd0;
    assign rom_im[67] = 9'sd0;
    assign rom_im[68] = 9'sd0;
    assign rom_im[69] = 9'sd0;
    assign rom_im[70] = 9'sd0;
    assign rom_im[71] = 9'sd0;
    assign rom_im[72] = 9'sd0;
    assign rom_im[73] = 9'sd0;
    assign rom_im[74] = 9'sd0;
    assign rom_im[75] = 9'sd0;
    assign rom_im[76] = 9'sd0;
    assign rom_im[77] = 9'sd0;
    assign rom_im[78] = 9'sd0;
    assign rom_im[79] = 9'sd0;
    assign rom_im[80] = 9'sd0;
    assign rom_im[81] = 9'sd0;
    assign rom_im[82] = 9'sd0;
    assign rom_im[83] = 9'sd0;
    assign rom_im[84] = 9'sd0;
    assign rom_im[85] = 9'sd0;
    assign rom_im[86] = 9'sd0;
    assign rom_im[87] = 9'sd0;
    assign rom_im[88] = 9'sd0;
    assign rom_im[89] = 9'sd0;
    assign rom_im[90] = 9'sd0;
    assign rom_im[91] = 9'sd0;
    assign rom_im[92] = 9'sd0;
    assign rom_im[93] = 9'sd0;
    assign rom_im[94] = 9'sd0;
    assign rom_im[95] = 9'sd0;
    assign rom_im[96] = 9'sd0;
    assign rom_im[97] = 9'sd0;
    assign rom_im[98] = 9'sd0;
    assign rom_im[99] = 9'sd0;
    assign rom_im[100] = 9'sd0;
    assign rom_im[101] = 9'sd0;
    assign rom_im[102] = 9'sd0;
    assign rom_im[103] = 9'sd0;
    assign rom_im[104] = 9'sd0;
    assign rom_im[105] = 9'sd0;
    assign rom_im[106] = 9'sd0;
    assign rom_im[107] = 9'sd0;
    assign rom_im[108] = 9'sd0;
    assign rom_im[109] = 9'sd0;
    assign rom_im[110] = 9'sd0;
    assign rom_im[111] = 9'sd0;
    assign rom_im[112] = 9'sd0;
    assign rom_im[113] = 9'sd0;
    assign rom_im[114] = 9'sd0;
    assign rom_im[115] = 9'sd0;
    assign rom_im[116] = 9'sd0;
    assign rom_im[117] = 9'sd0;
    assign rom_im[118] = 9'sd0;
    assign rom_im[119] = 9'sd0;
    assign rom_im[120] = 9'sd0;
    assign rom_im[121] = 9'sd0;
    assign rom_im[122] = 9'sd0;
    assign rom_im[123] = 9'sd0;
    assign rom_im[124] = 9'sd0;
    assign rom_im[125] = 9'sd0;
    assign rom_im[126] = 9'sd0;
    assign rom_im[127] = 9'sd0;
    assign rom_im[128] = 9'sd0;
    assign rom_im[129] = 9'sd0;
    assign rom_im[130] = 9'sd0;
    assign rom_im[131] = 9'sd0;
    assign rom_im[132] = 9'sd0;
    assign rom_im[133] = 9'sd0;
    assign rom_im[134] = 9'sd0;
    assign rom_im[135] = 9'sd0;
    assign rom_im[136] = 9'sd0;
    assign rom_im[137] = 9'sd0;
    assign rom_im[138] = 9'sd0;
    assign rom_im[139] = 9'sd0;
    assign rom_im[140] = 9'sd0;
    assign rom_im[141] = 9'sd0;
    assign rom_im[142] = 9'sd0;
    assign rom_im[143] = 9'sd0;
    assign rom_im[144] = 9'sd0;
    assign rom_im[145] = 9'sd0;
    assign rom_im[146] = 9'sd0;
    assign rom_im[147] = 9'sd0;
    assign rom_im[148] = 9'sd0;
    assign rom_im[149] = 9'sd0;
    assign rom_im[150] = 9'sd0;
    assign rom_im[151] = 9'sd0;
    assign rom_im[152] = 9'sd0;
    assign rom_im[153] = 9'sd0;
    assign rom_im[154] = 9'sd0;
    assign rom_im[155] = 9'sd0;
    assign rom_im[156] = 9'sd0;
    assign rom_im[157] = 9'sd0;
    assign rom_im[158] = 9'sd0;
    assign rom_im[159] = 9'sd0;
    assign rom_im[160] = 9'sd0;
    assign rom_im[161] = 9'sd0;
    assign rom_im[162] = 9'sd0;
    assign rom_im[163] = 9'sd0;
    assign rom_im[164] = 9'sd0;
    assign rom_im[165] = 9'sd0;
    assign rom_im[166] = 9'sd0;
    assign rom_im[167] = 9'sd0;
    assign rom_im[168] = 9'sd0;
    assign rom_im[169] = 9'sd0;
    assign rom_im[170] = 9'sd0;
    assign rom_im[171] = 9'sd0;
    assign rom_im[172] = 9'sd0;
    assign rom_im[173] = 9'sd0;
    assign rom_im[174] = 9'sd0;
    assign rom_im[175] = 9'sd0;
    assign rom_im[176] = 9'sd0;
    assign rom_im[177] = 9'sd0;
    assign rom_im[178] = 9'sd0;
    assign rom_im[179] = 9'sd0;
    assign rom_im[180] = 9'sd0;
    assign rom_im[181] = 9'sd0;
    assign rom_im[182] = 9'sd0;
    assign rom_im[183] = 9'sd0;
    assign rom_im[184] = 9'sd0;
    assign rom_im[185] = 9'sd0;
    assign rom_im[186] = 9'sd0;
    assign rom_im[187] = 9'sd0;
    assign rom_im[188] = 9'sd0;
    assign rom_im[189] = 9'sd0;
    assign rom_im[190] = 9'sd0;
    assign rom_im[191] = 9'sd0;
    assign rom_im[192] = 9'sd0;
    assign rom_im[193] = 9'sd0;
    assign rom_im[194] = 9'sd0;
    assign rom_im[195] = 9'sd0;
    assign rom_im[196] = 9'sd0;
    assign rom_im[197] = 9'sd0;
    assign rom_im[198] = 9'sd0;
    assign rom_im[199] = 9'sd0;
    assign rom_im[200] = 9'sd0;
    assign rom_im[201] = 9'sd0;
    assign rom_im[202] = 9'sd0;
    assign rom_im[203] = 9'sd0;
    assign rom_im[204] = 9'sd0;
    assign rom_im[205] = 9'sd0;
    assign rom_im[206] = 9'sd0;
    assign rom_im[207] = 9'sd0;
    assign rom_im[208] = 9'sd0;
    assign rom_im[209] = 9'sd0;
    assign rom_im[210] = 9'sd0;
    assign rom_im[211] = 9'sd0;
    assign rom_im[212] = 9'sd0;
    assign rom_im[213] = 9'sd0;
    assign rom_im[214] = 9'sd0;
    assign rom_im[215] = 9'sd0;
    assign rom_im[216] = 9'sd0;
    assign rom_im[217] = 9'sd0;
    assign rom_im[218] = 9'sd0;
    assign rom_im[219] = 9'sd0;
    assign rom_im[220] = 9'sd0;
    assign rom_im[221] = 9'sd0;
    assign rom_im[222] = 9'sd0;
    assign rom_im[223] = 9'sd0;
    assign rom_im[224] = 9'sd0;
    assign rom_im[225] = 9'sd0;
    assign rom_im[226] = 9'sd0;
    assign rom_im[227] = 9'sd0;
    assign rom_im[228] = 9'sd0;
    assign rom_im[229] = 9'sd0;
    assign rom_im[230] = 9'sd0;
    assign rom_im[231] = 9'sd0;
    assign rom_im[232] = 9'sd0;
    assign rom_im[233] = 9'sd0;
    assign rom_im[234] = 9'sd0;
    assign rom_im[235] = 9'sd0;
    assign rom_im[236] = 9'sd0;
    assign rom_im[237] = 9'sd0;
    assign rom_im[238] = 9'sd0;
    assign rom_im[239] = 9'sd0;
    assign rom_im[240] = 9'sd0;
    assign rom_im[241] = 9'sd0;
    assign rom_im[242] = 9'sd0;
    assign rom_im[243] = 9'sd0;
    assign rom_im[244] = 9'sd0;
    assign rom_im[245] = 9'sd0;
    assign rom_im[246] = 9'sd0;
    assign rom_im[247] = 9'sd0;
    assign rom_im[248] = 9'sd0;
    assign rom_im[249] = 9'sd0;
    assign rom_im[250] = 9'sd0;
    assign rom_im[251] = 9'sd0;
    assign rom_im[252] = 9'sd0;
    assign rom_im[253] = 9'sd0;
    assign rom_im[254] = 9'sd0;
    assign rom_im[255] = 9'sd0;
    assign rom_im[256] = 9'sd0;
    assign rom_im[257] = 9'sd0;
    assign rom_im[258] = 9'sd0;
    assign rom_im[259] = 9'sd0;
    assign rom_im[260] = 9'sd0;
    assign rom_im[261] = 9'sd0;
    assign rom_im[262] = 9'sd0;
    assign rom_im[263] = 9'sd0;
    assign rom_im[264] = 9'sd0;
    assign rom_im[265] = 9'sd0;
    assign rom_im[266] = 9'sd0;
    assign rom_im[267] = 9'sd0;
    assign rom_im[268] = 9'sd0;
    assign rom_im[269] = 9'sd0;
    assign rom_im[270] = 9'sd0;
    assign rom_im[271] = 9'sd0;
    assign rom_im[272] = 9'sd0;
    assign rom_im[273] = 9'sd0;
    assign rom_im[274] = 9'sd0;
    assign rom_im[275] = 9'sd0;
    assign rom_im[276] = 9'sd0;
    assign rom_im[277] = 9'sd0;
    assign rom_im[278] = 9'sd0;
    assign rom_im[279] = 9'sd0;
    assign rom_im[280] = 9'sd0;
    assign rom_im[281] = 9'sd0;
    assign rom_im[282] = 9'sd0;
    assign rom_im[283] = 9'sd0;
    assign rom_im[284] = 9'sd0;
    assign rom_im[285] = 9'sd0;
    assign rom_im[286] = 9'sd0;
    assign rom_im[287] = 9'sd0;
    assign rom_im[288] = 9'sd0;
    assign rom_im[289] = 9'sd0;
    assign rom_im[290] = 9'sd0;
    assign rom_im[291] = 9'sd0;
    assign rom_im[292] = 9'sd0;
    assign rom_im[293] = 9'sd0;
    assign rom_im[294] = 9'sd0;
    assign rom_im[295] = 9'sd0;
    assign rom_im[296] = 9'sd0;
    assign rom_im[297] = 9'sd0;
    assign rom_im[298] = 9'sd0;
    assign rom_im[299] = 9'sd0;
    assign rom_im[300] = 9'sd0;
    assign rom_im[301] = 9'sd0;
    assign rom_im[302] = 9'sd0;
    assign rom_im[303] = 9'sd0;
    assign rom_im[304] = 9'sd0;
    assign rom_im[305] = 9'sd0;
    assign rom_im[306] = 9'sd0;
    assign rom_im[307] = 9'sd0;
    assign rom_im[308] = 9'sd0;
    assign rom_im[309] = 9'sd0;
    assign rom_im[310] = 9'sd0;
    assign rom_im[311] = 9'sd0;
    assign rom_im[312] = 9'sd0;
    assign rom_im[313] = 9'sd0;
    assign rom_im[314] = 9'sd0;
    assign rom_im[315] = 9'sd0;
    assign rom_im[316] = 9'sd0;
    assign rom_im[317] = 9'sd0;
    assign rom_im[318] = 9'sd0;
    assign rom_im[319] = 9'sd0;
    assign rom_im[320] = 9'sd0;
    assign rom_im[321] = 9'sd0;
    assign rom_im[322] = 9'sd0;
    assign rom_im[323] = 9'sd0;
    assign rom_im[324] = 9'sd0;
    assign rom_im[325] = 9'sd0;
    assign rom_im[326] = 9'sd0;
    assign rom_im[327] = 9'sd0;
    assign rom_im[328] = 9'sd0;
    assign rom_im[329] = 9'sd0;
    assign rom_im[330] = 9'sd0;
    assign rom_im[331] = 9'sd0;
    assign rom_im[332] = 9'sd0;
    assign rom_im[333] = 9'sd0;
    assign rom_im[334] = 9'sd0;
    assign rom_im[335] = 9'sd0;
    assign rom_im[336] = 9'sd0;
    assign rom_im[337] = 9'sd0;
    assign rom_im[338] = 9'sd0;
    assign rom_im[339] = 9'sd0;
    assign rom_im[340] = 9'sd0;
    assign rom_im[341] = 9'sd0;
    assign rom_im[342] = 9'sd0;
    assign rom_im[343] = 9'sd0;
    assign rom_im[344] = 9'sd0;
    assign rom_im[345] = 9'sd0;
    assign rom_im[346] = 9'sd0;
    assign rom_im[347] = 9'sd0;
    assign rom_im[348] = 9'sd0;
    assign rom_im[349] = 9'sd0;
    assign rom_im[350] = 9'sd0;
    assign rom_im[351] = 9'sd0;
    assign rom_im[352] = 9'sd0;
    assign rom_im[353] = 9'sd0;
    assign rom_im[354] = 9'sd0;
    assign rom_im[355] = 9'sd0;
    assign rom_im[356] = 9'sd0;
    assign rom_im[357] = 9'sd0;
    assign rom_im[358] = 9'sd0;
    assign rom_im[359] = 9'sd0;
    assign rom_im[360] = 9'sd0;
    assign rom_im[361] = 9'sd0;
    assign rom_im[362] = 9'sd0;
    assign rom_im[363] = 9'sd0;
    assign rom_im[364] = 9'sd0;
    assign rom_im[365] = 9'sd0;
    assign rom_im[366] = 9'sd0;
    assign rom_im[367] = 9'sd0;
    assign rom_im[368] = 9'sd0;
    assign rom_im[369] = 9'sd0;
    assign rom_im[370] = 9'sd0;
    assign rom_im[371] = 9'sd0;
    assign rom_im[372] = 9'sd0;
    assign rom_im[373] = 9'sd0;
    assign rom_im[374] = 9'sd0;
    assign rom_im[375] = 9'sd0;
    assign rom_im[376] = 9'sd0;
    assign rom_im[377] = 9'sd0;
    assign rom_im[378] = 9'sd0;
    assign rom_im[379] = 9'sd0;
    assign rom_im[380] = 9'sd0;
    assign rom_im[381] = 9'sd0;
    assign rom_im[382] = 9'sd0;
    assign rom_im[383] = 9'sd0;
    assign rom_im[384] = 9'sd0;
    assign rom_im[385] = 9'sd0;
    assign rom_im[386] = 9'sd0;
    assign rom_im[387] = 9'sd0;
    assign rom_im[388] = 9'sd0;
    assign rom_im[389] = 9'sd0;
    assign rom_im[390] = 9'sd0;
    assign rom_im[391] = 9'sd0;
    assign rom_im[392] = 9'sd0;
    assign rom_im[393] = 9'sd0;
    assign rom_im[394] = 9'sd0;
    assign rom_im[395] = 9'sd0;
    assign rom_im[396] = 9'sd0;
    assign rom_im[397] = 9'sd0;
    assign rom_im[398] = 9'sd0;
    assign rom_im[399] = 9'sd0;
    assign rom_im[400] = 9'sd0;
    assign rom_im[401] = 9'sd0;
    assign rom_im[402] = 9'sd0;
    assign rom_im[403] = 9'sd0;
    assign rom_im[404] = 9'sd0;
    assign rom_im[405] = 9'sd0;
    assign rom_im[406] = 9'sd0;
    assign rom_im[407] = 9'sd0;
    assign rom_im[408] = 9'sd0;
    assign rom_im[409] = 9'sd0;
    assign rom_im[410] = 9'sd0;
    assign rom_im[411] = 9'sd0;
    assign rom_im[412] = 9'sd0;
    assign rom_im[413] = 9'sd0;
    assign rom_im[414] = 9'sd0;
    assign rom_im[415] = 9'sd0;
    assign rom_im[416] = 9'sd0;
    assign rom_im[417] = 9'sd0;
    assign rom_im[418] = 9'sd0;
    assign rom_im[419] = 9'sd0;
    assign rom_im[420] = 9'sd0;
    assign rom_im[421] = 9'sd0;
    assign rom_im[422] = 9'sd0;
    assign rom_im[423] = 9'sd0;
    assign rom_im[424] = 9'sd0;
    assign rom_im[425] = 9'sd0;
    assign rom_im[426] = 9'sd0;
    assign rom_im[427] = 9'sd0;
    assign rom_im[428] = 9'sd0;
    assign rom_im[429] = 9'sd0;
    assign rom_im[430] = 9'sd0;
    assign rom_im[431] = 9'sd0;
    assign rom_im[432] = 9'sd0;
    assign rom_im[433] = 9'sd0;
    assign rom_im[434] = 9'sd0;
    assign rom_im[435] = 9'sd0;
    assign rom_im[436] = 9'sd0;
    assign rom_im[437] = 9'sd0;
    assign rom_im[438] = 9'sd0;
    assign rom_im[439] = 9'sd0;
    assign rom_im[440] = 9'sd0;
    assign rom_im[441] = 9'sd0;
    assign rom_im[442] = 9'sd0;
    assign rom_im[443] = 9'sd0;
    assign rom_im[444] = 9'sd0;
    assign rom_im[445] = 9'sd0;
    assign rom_im[446] = 9'sd0;
    assign rom_im[447] = 9'sd0;
    assign rom_im[448] = 9'sd0;
    assign rom_im[449] = 9'sd0;
    assign rom_im[450] = 9'sd0;
    assign rom_im[451] = 9'sd0;
    assign rom_im[452] = 9'sd0;
    assign rom_im[453] = 9'sd0;
    assign rom_im[454] = 9'sd0;
    assign rom_im[455] = 9'sd0;
    assign rom_im[456] = 9'sd0;
    assign rom_im[457] = 9'sd0;
    assign rom_im[458] = 9'sd0;
    assign rom_im[459] = 9'sd0;
    assign rom_im[460] = 9'sd0;
    assign rom_im[461] = 9'sd0;
    assign rom_im[462] = 9'sd0;
    assign rom_im[463] = 9'sd0;
    assign rom_im[464] = 9'sd0;
    assign rom_im[465] = 9'sd0;
    assign rom_im[466] = 9'sd0;
    assign rom_im[467] = 9'sd0;
    assign rom_im[468] = 9'sd0;
    assign rom_im[469] = 9'sd0;
    assign rom_im[470] = 9'sd0;
    assign rom_im[471] = 9'sd0;
    assign rom_im[472] = 9'sd0;
    assign rom_im[473] = 9'sd0;
    assign rom_im[474] = 9'sd0;
    assign rom_im[475] = 9'sd0;
    assign rom_im[476] = 9'sd0;
    assign rom_im[477] = 9'sd0;
    assign rom_im[478] = 9'sd0;
    assign rom_im[479] = 9'sd0;
    assign rom_im[480] = 9'sd0;
    assign rom_im[481] = 9'sd0;
    assign rom_im[482] = 9'sd0;
    assign rom_im[483] = 9'sd0;
    assign rom_im[484] = 9'sd0;
    assign rom_im[485] = 9'sd0;
    assign rom_im[486] = 9'sd0;
    assign rom_im[487] = 9'sd0;
    assign rom_im[488] = 9'sd0;
    assign rom_im[489] = 9'sd0;
    assign rom_im[490] = 9'sd0;
    assign rom_im[491] = 9'sd0;
    assign rom_im[492] = 9'sd0;
    assign rom_im[493] = 9'sd0;
    assign rom_im[494] = 9'sd0;
    assign rom_im[495] = 9'sd0;
    assign rom_im[496] = 9'sd0;
    assign rom_im[497] = 9'sd0;
    assign rom_im[498] = 9'sd0;
    assign rom_im[499] = 9'sd0;
    assign rom_im[500] = 9'sd0;
    assign rom_im[501] = 9'sd0;
    assign rom_im[502] = 9'sd0;
    assign rom_im[503] = 9'sd0;
    assign rom_im[504] = 9'sd0;
    assign rom_im[505] = 9'sd0;
    assign rom_im[506] = 9'sd0;
    assign rom_im[507] = 9'sd0;
    assign rom_im[508] = 9'sd0;
    assign rom_im[509] = 9'sd0;
    assign rom_im[510] = 9'sd0;
    assign rom_im[511] = 9'sd0;

    // cos_rom_i_assign.txt
    assign rom_re[0] = 9'sd63;
    assign rom_re[1] = 9'sd64;
    assign rom_re[2] = 9'sd64;
    assign rom_re[3] = 9'sd64;
    assign rom_re[4] = 9'sd64;
    assign rom_re[5] = 9'sd64;
    assign rom_re[6] = 9'sd64;
    assign rom_re[7] = 9'sd64;
    assign rom_re[8] = 9'sd64;
    assign rom_re[9] = 9'sd64;
    assign rom_re[10] = 9'sd64;
    assign rom_re[11] = 9'sd63;
    assign rom_re[12] = 9'sd63;
    assign rom_re[13] = 9'sd63;
    assign rom_re[14] = 9'sd63;
    assign rom_re[15] = 9'sd63;
    assign rom_re[16] = 9'sd63;
    assign rom_re[17] = 9'sd63;
    assign rom_re[18] = 9'sd62;
    assign rom_re[19] = 9'sd62;
    assign rom_re[20] = 9'sd62;
    assign rom_re[21] = 9'sd62;
    assign rom_re[22] = 9'sd62;
    assign rom_re[23] = 9'sd61;
    assign rom_re[24] = 9'sd61;
    assign rom_re[25] = 9'sd61;
    assign rom_re[26] = 9'sd61;
    assign rom_re[27] = 9'sd61;
    assign rom_re[28] = 9'sd60;
    assign rom_re[29] = 9'sd60;
    assign rom_re[30] = 9'sd60;
    assign rom_re[31] = 9'sd59;
    assign rom_re[32] = 9'sd59;
    assign rom_re[33] = 9'sd59;
    assign rom_re[34] = 9'sd59;
    assign rom_re[35] = 9'sd58;
    assign rom_re[36] = 9'sd58;
    assign rom_re[37] = 9'sd58;
    assign rom_re[38] = 9'sd57;
    assign rom_re[39] = 9'sd57;
    assign rom_re[40] = 9'sd56;
    assign rom_re[41] = 9'sd56;
    assign rom_re[42] = 9'sd56;
    assign rom_re[43] = 9'sd55;
    assign rom_re[44] = 9'sd55;
    assign rom_re[45] = 9'sd54;
    assign rom_re[46] = 9'sd54;
    assign rom_re[47] = 9'sd54;
    assign rom_re[48] = 9'sd53;
    assign rom_re[49] = 9'sd53;
    assign rom_re[50] = 9'sd52;
    assign rom_re[51] = 9'sd52;
    assign rom_re[52] = 9'sd51;
    assign rom_re[53] = 9'sd51;
    assign rom_re[54] = 9'sd50;
    assign rom_re[55] = 9'sd50;
    assign rom_re[56] = 9'sd49;
    assign rom_re[57] = 9'sd49;
    assign rom_re[58] = 9'sd48;
    assign rom_re[59] = 9'sd48;
    assign rom_re[60] = 9'sd47;
    assign rom_re[61] = 9'sd47;
    assign rom_re[62] = 9'sd46;
    assign rom_re[63] = 9'sd46;
    assign rom_re[64] = 9'sd45;
    assign rom_re[65] = 9'sd45;
    assign rom_re[66] = 9'sd44;
    assign rom_re[67] = 9'sd44;
    assign rom_re[68] = 9'sd43;
    assign rom_re[69] = 9'sd42;
    assign rom_re[70] = 9'sd42;
    assign rom_re[71] = 9'sd41;
    assign rom_re[72] = 9'sd41;
    assign rom_re[73] = 9'sd40;
    assign rom_re[74] = 9'sd39;
    assign rom_re[75] = 9'sd39;
    assign rom_re[76] = 9'sd38;
    assign rom_re[77] = 9'sd37;
    assign rom_re[78] = 9'sd37;
    assign rom_re[79] = 9'sd36;
    assign rom_re[80] = 9'sd36;
    assign rom_re[81] = 9'sd35;
    assign rom_re[82] = 9'sd34;
    assign rom_re[83] = 9'sd34;
    assign rom_re[84] = 9'sd33;
    assign rom_re[85] = 9'sd32;
    assign rom_re[86] = 9'sd32;
    assign rom_re[87] = 9'sd31;
    assign rom_re[88] = 9'sd30;
    assign rom_re[89] = 9'sd29;
    assign rom_re[90] = 9'sd29;
    assign rom_re[91] = 9'sd28;
    assign rom_re[92] = 9'sd27;
    assign rom_re[93] = 9'sd27;
    assign rom_re[94] = 9'sd26;
    assign rom_re[95] = 9'sd25;
    assign rom_re[96] = 9'sd24;
    assign rom_re[97] = 9'sd24;
    assign rom_re[98] = 9'sd23;
    assign rom_re[99] = 9'sd22;
    assign rom_re[100] = 9'sd22;
    assign rom_re[101] = 9'sd21;
    assign rom_re[102] = 9'sd20;
    assign rom_re[103] = 9'sd19;
    assign rom_re[104] = 9'sd19;
    assign rom_re[105] = 9'sd18;
    assign rom_re[106] = 9'sd17;
    assign rom_re[107] = 9'sd16;
    assign rom_re[108] = 9'sd16;
    assign rom_re[109] = 9'sd15;
    assign rom_re[110] = 9'sd14;
    assign rom_re[111] = 9'sd13;
    assign rom_re[112] = 9'sd12;
    assign rom_re[113] = 9'sd12;
    assign rom_re[114] = 9'sd11;
    assign rom_re[115] = 9'sd10;
    assign rom_re[116] = 9'sd9;
    assign rom_re[117] = 9'sd9;
    assign rom_re[118] = 9'sd8;
    assign rom_re[119] = 9'sd7;
    assign rom_re[120] = 9'sd6;
    assign rom_re[121] = 9'sd5;
    assign rom_re[122] = 9'sd5;
    assign rom_re[123] = 9'sd4;
    assign rom_re[124] = 9'sd3;
    assign rom_re[125] = 9'sd2;
    assign rom_re[126] = 9'sd2;
    assign rom_re[127] = 9'sd1;
    assign rom_re[128] = 9'sd0;
    assign rom_re[129] = -9'sd1;
    assign rom_re[130] = -9'sd2;
    assign rom_re[131] = -9'sd2;
    assign rom_re[132] = -9'sd3;
    assign rom_re[133] = -9'sd4;
    assign rom_re[134] = -9'sd5;
    assign rom_re[135] = -9'sd5;
    assign rom_re[136] = -9'sd6;
    assign rom_re[137] = -9'sd7;
    assign rom_re[138] = -9'sd8;
    assign rom_re[139] = -9'sd9;
    assign rom_re[140] = -9'sd9;
    assign rom_re[141] = -9'sd10;
    assign rom_re[142] = -9'sd11;
    assign rom_re[143] = -9'sd12;
    assign rom_re[144] = -9'sd12;
    assign rom_re[145] = -9'sd13;
    assign rom_re[146] = -9'sd14;
    assign rom_re[147] = -9'sd15;
    assign rom_re[148] = -9'sd16;
    assign rom_re[149] = -9'sd16;
    assign rom_re[150] = -9'sd17;
    assign rom_re[151] = -9'sd18;
    assign rom_re[152] = -9'sd19;
    assign rom_re[153] = -9'sd19;
    assign rom_re[154] = -9'sd20;
    assign rom_re[155] = -9'sd21;
    assign rom_re[156] = -9'sd22;
    assign rom_re[157] = -9'sd22;
    assign rom_re[158] = -9'sd23;
    assign rom_re[159] = -9'sd24;
    assign rom_re[160] = -9'sd24;
    assign rom_re[161] = -9'sd25;
    assign rom_re[162] = -9'sd26;
    assign rom_re[163] = -9'sd27;
    assign rom_re[164] = -9'sd27;
    assign rom_re[165] = -9'sd28;
    assign rom_re[166] = -9'sd29;
    assign rom_re[167] = -9'sd29;
    assign rom_re[168] = -9'sd30;
    assign rom_re[169] = -9'sd31;
    assign rom_re[170] = -9'sd32;
    assign rom_re[171] = -9'sd32;
    assign rom_re[172] = -9'sd33;
    assign rom_re[173] = -9'sd34;
    assign rom_re[174] = -9'sd34;
    assign rom_re[175] = -9'sd35;
    assign rom_re[176] = -9'sd36;
    assign rom_re[177] = -9'sd36;
    assign rom_re[178] = -9'sd37;
    assign rom_re[179] = -9'sd37;
    assign rom_re[180] = -9'sd38;
    assign rom_re[181] = -9'sd39;
    assign rom_re[182] = -9'sd39;
    assign rom_re[183] = -9'sd40;
    assign rom_re[184] = -9'sd41;
    assign rom_re[185] = -9'sd41;
    assign rom_re[186] = -9'sd42;
    assign rom_re[187] = -9'sd42;
    assign rom_re[188] = -9'sd43;
    assign rom_re[189] = -9'sd44;
    assign rom_re[190] = -9'sd44;
    assign rom_re[191] = -9'sd45;
    assign rom_re[192] = -9'sd45;
    assign rom_re[193] = -9'sd46;
    assign rom_re[194] = -9'sd46;
    assign rom_re[195] = -9'sd47;
    assign rom_re[196] = -9'sd47;
    assign rom_re[197] = -9'sd48;
    assign rom_re[198] = -9'sd48;
    assign rom_re[199] = -9'sd49;
    assign rom_re[200] = -9'sd49;
    assign rom_re[201] = -9'sd50;
    assign rom_re[202] = -9'sd50;
    assign rom_re[203] = -9'sd51;
    assign rom_re[204] = -9'sd51;
    assign rom_re[205] = -9'sd52;
    assign rom_re[206] = -9'sd52;
    assign rom_re[207] = -9'sd53;
    assign rom_re[208] = -9'sd53;
    assign rom_re[209] = -9'sd54;
    assign rom_re[210] = -9'sd54;
    assign rom_re[211] = -9'sd54;
    assign rom_re[212] = -9'sd55;
    assign rom_re[213] = -9'sd55;
    assign rom_re[214] = -9'sd56;
    assign rom_re[215] = -9'sd56;
    assign rom_re[216] = -9'sd56;
    assign rom_re[217] = -9'sd57;
    assign rom_re[218] = -9'sd57;
    assign rom_re[219] = -9'sd58;
    assign rom_re[220] = -9'sd58;
    assign rom_re[221] = -9'sd58;
    assign rom_re[222] = -9'sd59;
    assign rom_re[223] = -9'sd59;
    assign rom_re[224] = -9'sd59;
    assign rom_re[225] = -9'sd59;
    assign rom_re[226] = -9'sd60;
    assign rom_re[227] = -9'sd60;
    assign rom_re[228] = -9'sd60;
    assign rom_re[229] = -9'sd61;
    assign rom_re[230] = -9'sd61;
    assign rom_re[231] = -9'sd61;
    assign rom_re[232] = -9'sd61;
    assign rom_re[233] = -9'sd61;
    assign rom_re[234] = -9'sd62;
    assign rom_re[235] = -9'sd62;
    assign rom_re[236] = -9'sd62;
    assign rom_re[237] = -9'sd62;
    assign rom_re[238] = -9'sd62;
    assign rom_re[239] = -9'sd63;
    assign rom_re[240] = -9'sd63;
    assign rom_re[241] = -9'sd63;
    assign rom_re[242] = -9'sd63;
    assign rom_re[243] = -9'sd63;
    assign rom_re[244] = -9'sd63;
    assign rom_re[245] = -9'sd63;
    assign rom_re[246] = -9'sd64;
    assign rom_re[247] = -9'sd64;
    assign rom_re[248] = -9'sd64;
    assign rom_re[249] = -9'sd64;
    assign rom_re[250] = -9'sd64;
    assign rom_re[251] = -9'sd64;
    assign rom_re[252] = -9'sd64;
    assign rom_re[253] = -9'sd64;
    assign rom_re[254] = -9'sd64;
    assign rom_re[255] = -9'sd64;
    assign rom_re[256] = -9'sd64;
    assign rom_re[257] = -9'sd64;
    assign rom_re[258] = -9'sd64;
    assign rom_re[259] = -9'sd64;
    assign rom_re[260] = -9'sd64;
    assign rom_re[261] = -9'sd64;
    assign rom_re[262] = -9'sd64;
    assign rom_re[263] = -9'sd64;
    assign rom_re[264] = -9'sd64;
    assign rom_re[265] = -9'sd64;
    assign rom_re[266] = -9'sd64;
    assign rom_re[267] = -9'sd63;
    assign rom_re[268] = -9'sd63;
    assign rom_re[269] = -9'sd63;
    assign rom_re[270] = -9'sd63;
    assign rom_re[271] = -9'sd63;
    assign rom_re[272] = -9'sd63;
    assign rom_re[273] = -9'sd63;
    assign rom_re[274] = -9'sd62;
    assign rom_re[275] = -9'sd62;
    assign rom_re[276] = -9'sd62;
    assign rom_re[277] = -9'sd62;
    assign rom_re[278] = -9'sd62;
    assign rom_re[279] = -9'sd61;
    assign rom_re[280] = -9'sd61;
    assign rom_re[281] = -9'sd61;
    assign rom_re[282] = -9'sd61;
    assign rom_re[283] = -9'sd61;
    assign rom_re[284] = -9'sd60;
    assign rom_re[285] = -9'sd60;
    assign rom_re[286] = -9'sd60;
    assign rom_re[287] = -9'sd59;
    assign rom_re[288] = -9'sd59;
    assign rom_re[289] = -9'sd59;
    assign rom_re[290] = -9'sd59;
    assign rom_re[291] = -9'sd58;
    assign rom_re[292] = -9'sd58;
    assign rom_re[293] = -9'sd58;
    assign rom_re[294] = -9'sd57;
    assign rom_re[295] = -9'sd57;
    assign rom_re[296] = -9'sd56;
    assign rom_re[297] = -9'sd56;
    assign rom_re[298] = -9'sd56;
    assign rom_re[299] = -9'sd55;
    assign rom_re[300] = -9'sd55;
    assign rom_re[301] = -9'sd54;
    assign rom_re[302] = -9'sd54;
    assign rom_re[303] = -9'sd54;
    assign rom_re[304] = -9'sd53;
    assign rom_re[305] = -9'sd53;
    assign rom_re[306] = -9'sd52;
    assign rom_re[307] = -9'sd52;
    assign rom_re[308] = -9'sd51;
    assign rom_re[309] = -9'sd51;
    assign rom_re[310] = -9'sd50;
    assign rom_re[311] = -9'sd50;
    assign rom_re[312] = -9'sd49;
    assign rom_re[313] = -9'sd49;
    assign rom_re[314] = -9'sd48;
    assign rom_re[315] = -9'sd48;
    assign rom_re[316] = -9'sd47;
    assign rom_re[317] = -9'sd47;
    assign rom_re[318] = -9'sd46;
    assign rom_re[319] = -9'sd46;
    assign rom_re[320] = -9'sd45;
    assign rom_re[321] = -9'sd45;
    assign rom_re[322] = -9'sd44;
    assign rom_re[323] = -9'sd44;
    assign rom_re[324] = -9'sd43;
    assign rom_re[325] = -9'sd42;
    assign rom_re[326] = -9'sd42;
    assign rom_re[327] = -9'sd41;
    assign rom_re[328] = -9'sd41;
    assign rom_re[329] = -9'sd40;
    assign rom_re[330] = -9'sd39;
    assign rom_re[331] = -9'sd39;
    assign rom_re[332] = -9'sd38;
    assign rom_re[333] = -9'sd37;
    assign rom_re[334] = -9'sd37;
    assign rom_re[335] = -9'sd36;
    assign rom_re[336] = -9'sd36;
    assign rom_re[337] = -9'sd35;
    assign rom_re[338] = -9'sd34;
    assign rom_re[339] = -9'sd34;
    assign rom_re[340] = -9'sd33;
    assign rom_re[341] = -9'sd32;
    assign rom_re[342] = -9'sd32;
    assign rom_re[343] = -9'sd31;
    assign rom_re[344] = -9'sd30;
    assign rom_re[345] = -9'sd29;
    assign rom_re[346] = -9'sd29;
    assign rom_re[347] = -9'sd28;
    assign rom_re[348] = -9'sd27;
    assign rom_re[349] = -9'sd27;
    assign rom_re[350] = -9'sd26;
    assign rom_re[351] = -9'sd25;
    assign rom_re[352] = -9'sd24;
    assign rom_re[353] = -9'sd24;
    assign rom_re[354] = -9'sd23;
    assign rom_re[355] = -9'sd22;
    assign rom_re[356] = -9'sd22;
    assign rom_re[357] = -9'sd21;
    assign rom_re[358] = -9'sd20;
    assign rom_re[359] = -9'sd19;
    assign rom_re[360] = -9'sd19;
    assign rom_re[361] = -9'sd18;
    assign rom_re[362] = -9'sd17;
    assign rom_re[363] = -9'sd16;
    assign rom_re[364] = -9'sd16;
    assign rom_re[365] = -9'sd15;
    assign rom_re[366] = -9'sd14;
    assign rom_re[367] = -9'sd13;
    assign rom_re[368] = -9'sd12;
    assign rom_re[369] = -9'sd12;
    assign rom_re[370] = -9'sd11;
    assign rom_re[371] = -9'sd10;
    assign rom_re[372] = -9'sd9;
    assign rom_re[373] = -9'sd9;
    assign rom_re[374] = -9'sd8;
    assign rom_re[375] = -9'sd7;
    assign rom_re[376] = -9'sd6;
    assign rom_re[377] = -9'sd5;
    assign rom_re[378] = -9'sd5;
    assign rom_re[379] = -9'sd4;
    assign rom_re[380] = -9'sd3;
    assign rom_re[381] = -9'sd2;
    assign rom_re[382] = -9'sd2;
    assign rom_re[383] = -9'sd1;
    assign rom_re[384] = 9'sd0;
    assign rom_re[385] = 9'sd1;
    assign rom_re[386] = 9'sd2;
    assign rom_re[387] = 9'sd2;
    assign rom_re[388] = 9'sd3;
    assign rom_re[389] = 9'sd4;
    assign rom_re[390] = 9'sd5;
    assign rom_re[391] = 9'sd5;
    assign rom_re[392] = 9'sd6;
    assign rom_re[393] = 9'sd7;
    assign rom_re[394] = 9'sd8;
    assign rom_re[395] = 9'sd9;
    assign rom_re[396] = 9'sd9;
    assign rom_re[397] = 9'sd10;
    assign rom_re[398] = 9'sd11;
    assign rom_re[399] = 9'sd12;
    assign rom_re[400] = 9'sd12;
    assign rom_re[401] = 9'sd13;
    assign rom_re[402] = 9'sd14;
    assign rom_re[403] = 9'sd15;
    assign rom_re[404] = 9'sd16;
    assign rom_re[405] = 9'sd16;
    assign rom_re[406] = 9'sd17;
    assign rom_re[407] = 9'sd18;
    assign rom_re[408] = 9'sd19;
    assign rom_re[409] = 9'sd19;
    assign rom_re[410] = 9'sd20;
    assign rom_re[411] = 9'sd21;
    assign rom_re[412] = 9'sd22;
    assign rom_re[413] = 9'sd22;
    assign rom_re[414] = 9'sd23;
    assign rom_re[415] = 9'sd24;
    assign rom_re[416] = 9'sd24;
    assign rom_re[417] = 9'sd25;
    assign rom_re[418] = 9'sd26;
    assign rom_re[419] = 9'sd27;
    assign rom_re[420] = 9'sd27;
    assign rom_re[421] = 9'sd28;
    assign rom_re[422] = 9'sd29;
    assign rom_re[423] = 9'sd29;
    assign rom_re[424] = 9'sd30;
    assign rom_re[425] = 9'sd31;
    assign rom_re[426] = 9'sd32;
    assign rom_re[427] = 9'sd32;
    assign rom_re[428] = 9'sd33;
    assign rom_re[429] = 9'sd34;
    assign rom_re[430] = 9'sd34;
    assign rom_re[431] = 9'sd35;
    assign rom_re[432] = 9'sd36;
    assign rom_re[433] = 9'sd36;
    assign rom_re[434] = 9'sd37;
    assign rom_re[435] = 9'sd37;
    assign rom_re[436] = 9'sd38;
    assign rom_re[437] = 9'sd39;
    assign rom_re[438] = 9'sd39;
    assign rom_re[439] = 9'sd40;
    assign rom_re[440] = 9'sd41;
    assign rom_re[441] = 9'sd41;
    assign rom_re[442] = 9'sd42;
    assign rom_re[443] = 9'sd42;
    assign rom_re[444] = 9'sd43;
    assign rom_re[445] = 9'sd44;
    assign rom_re[446] = 9'sd44;
    assign rom_re[447] = 9'sd45;
    assign rom_re[448] = 9'sd45;
    assign rom_re[449] = 9'sd46;
    assign rom_re[450] = 9'sd46;
    assign rom_re[451] = 9'sd47;
    assign rom_re[452] = 9'sd47;
    assign rom_re[453] = 9'sd48;
    assign rom_re[454] = 9'sd48;
    assign rom_re[455] = 9'sd49;
    assign rom_re[456] = 9'sd49;
    assign rom_re[457] = 9'sd50;
    assign rom_re[458] = 9'sd50;
    assign rom_re[459] = 9'sd51;
    assign rom_re[460] = 9'sd51;
    assign rom_re[461] = 9'sd52;
    assign rom_re[462] = 9'sd52;
    assign rom_re[463] = 9'sd53;
    assign rom_re[464] = 9'sd53;
    assign rom_re[465] = 9'sd54;
    assign rom_re[466] = 9'sd54;
    assign rom_re[467] = 9'sd54;
    assign rom_re[468] = 9'sd55;
    assign rom_re[469] = 9'sd55;
    assign rom_re[470] = 9'sd56;
    assign rom_re[471] = 9'sd56;
    assign rom_re[472] = 9'sd56;
    assign rom_re[473] = 9'sd57;
    assign rom_re[474] = 9'sd57;
    assign rom_re[475] = 9'sd58;
    assign rom_re[476] = 9'sd58;
    assign rom_re[477] = 9'sd58;
    assign rom_re[478] = 9'sd59;
    assign rom_re[479] = 9'sd59;
    assign rom_re[480] = 9'sd59;
    assign rom_re[481] = 9'sd59;
    assign rom_re[482] = 9'sd60;
    assign rom_re[483] = 9'sd60;
    assign rom_re[484] = 9'sd60;
    assign rom_re[485] = 9'sd61;
    assign rom_re[486] = 9'sd61;
    assign rom_re[487] = 9'sd61;
    assign rom_re[488] = 9'sd61;
    assign rom_re[489] = 9'sd61;
    assign rom_re[490] = 9'sd62;
    assign rom_re[491] = 9'sd62;
    assign rom_re[492] = 9'sd62;
    assign rom_re[493] = 9'sd62;
    assign rom_re[494] = 9'sd62;
    assign rom_re[495] = 9'sd63;
    assign rom_re[496] = 9'sd63;
    assign rom_re[497] = 9'sd63;
    assign rom_re[498] = 9'sd63;
    assign rom_re[499] = 9'sd63;
    assign rom_re[500] = 9'sd63;
    assign rom_re[501] = 9'sd63;
    assign rom_re[502] = 9'sd64;
    assign rom_re[503] = 9'sd64;
    assign rom_re[504] = 9'sd64;
    assign rom_re[505] = 9'sd64;
    assign rom_re[506] = 9'sd64;
    assign rom_re[507] = 9'sd64;
    assign rom_re[508] = 9'sd64;
    assign rom_re[509] = 9'sd64;
    assign rom_re[510] = 9'sd64;
    assign rom_re[511] = 9'sd64;

endmodule




`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        $readmemh("code.mem", rom);
        /*
        //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _ op // R-Type
        rom[0] = 32'b0000000_00001_00010_000_00011_0110011; // add  x3, x1, x2   12 + 11 = 23
        rom[1] = 32'b0100000_00001_00010_000_00100_0110011; // sub  x4, x1, x2   12 - 11 = 1
        rom[2] = 32'b0000000_00100_00001_001_00101_0110011; // sll  x5, x4, x1   11 << 1 = 22
        rom[3] = 32'b0000000_00100_00101_101_00110_0110011; // srl  x6, x4, x5   22 >> 1 = 11
        rom[4] = 32'b0100000_00100_11111_101_00111_0110011; // sra  x7, x4, x31  -8 >>> 1 = -4 
        rom[5] = 32'b0000000_11111_00010_010_01000_0110011; // slt  x8, x2, x31   -8 < 1 ? = 1 
        rom[6] = 32'b0000000_11111_00010_011_01001_0110011; // sltu x9, x2, x31   u(-8) < 1 ? = 0
        rom[7] = 32'b0000000_00001_00010_100_01010_0110011; // xor  x10, x1, x2   11 ^ 12 = 7 (b0111)
        rom[8] = 32'b0000000_00001_00010_110_01011_0110011; // or   x11, x1, x2   11 | 12 = 15(b1111)
        rom[9] = 32'b0000000_00001_00010_111_01100_0110011; // and  x12, x1, x2   11 & 12 = 8(b1000)

        //rom[x]= 32'bimm12_imm[10:5]_rs2_rs1_f3_imm[4:1]_imm11_op // B-Type
        rom[10] = 32'b0_000000_00010_00010_000_0100_0_1100011;  // beq x2, x2, 8

        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
        rom[11] = 32'b0000000_00000_00000_000_00000_0000000;  // jump되서 생략됌.
        rom[12] = 32'b0000000_00001_00000_010_00100_0100011;  // sw x1, 4(x0)
        rom[13] = 32'b0000000_00001_00000_001_00110_0100011;  // sh x1, 6(x0)
        rom[14] = 32'b0000000_00001_00000_000_00101_0100011;  // sb x1, 5(x0)

        //rom[x]= 32'bimm12_imm[10:5]_rs2_rs1_f3_imm[4:1]_imm11_op // B-Type
        rom[15] = 32'b0_000000_00010_00010_001_0100_0_1100011;  // bne x2, x2, 8
        //rom[x]= 32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
        rom[16] = 32'b0000000_11111_00000_010_01000_0100011;  // sw x31, 8(x0)

        //rom[x]= 32'bimm12_imm[10:5]_rs2_rs1_f3_imm[4:1]_imm11_op // B-Type
        rom[17] = 32'b0_000000_00010_00001_110_0100_0_1100011;  // bltu x1, x2, 8
        rom[18] = 32'b0000000_00000_00000_000_00000_0000000;

        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
        rom[19] = 32'b000000001000_00000_000_00100_0000011;  // lb  x4, 6(x0)
        rom[20] = 32'b000000001000_00000_001_00101_0000011;  // lh  x5, 6(x0)
        rom[21] = 32'b000000001000_00000_010_00110_0000011;  // lw  x6, 8(x0)
        rom[22] = 32'b000000001000_00000_100_00111_0000011;  // lbu x7, 5(x0)
        rom[23] = 32'b000000001000_00000_101_01000_0000011;  // lhu x8, 8(x0)
        
        //rom[x]= 32'bimm12_imm[10:5]_rs2_rs1_f3_imm[4:1]_imm11_op // B-Type
        rom[24] = 32'b0_000000_00010_00001_111_0100_0_1100011;  // bgeu x1, x2, 8

        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type
        rom[25] = 32'b000000000100_00001_000_00100_0010011;  // addi  x4, x1, 4  11 + 4 = 15
        rom[26] = 32'b100000000000_00001_010_00101_0010011;  // slti  x5, x1, 12  11 < - = 1
        rom[27] = 32'b100000000000_00001_011_00110_0010011;  // sltiu x6, x1, 12  11 < + = 0
        rom[28] = 32'b000000000100_00001_100_00111_0010011;  // xori  x7, x1, 4  11 ^ 4 = 15
        rom[29] = 32'b000000010000_00001_110_01000_0010011;  // ori   x8, x1, 16 11 | 16 = 27
        rom[30] = 32'b000000000010_00001_111_01001_0010011;  // andi  x9, x1, 2 11 & 2 = 2
        rom[31] = 32'b000000000011_00001_001_01010_0010011;  // slli x10, x1, 1 // 32'b00001011 << 3
        rom[32] = 32'b000000000011_11110_101_01011_0010011;  // srli x11, x30, 1 // -32 >> 3
        rom[33] = 32'b010000000011_11110_101_01100_0010011;  // srai x12, x30, 1 // -32 >>> 3

        //rom[x]= 32'bimm12_imm[10:5]_rs2_rs1_f3_imm[4:1]_imm11_op // B-Type
        rom[34] = 32'b0_000000_00010_11110_100_0100_0_1100011;  // blt x30, x2, 8
        rom[35] = 32'b0000000_00000_00000_000_00000_0000000;
        rom[36] = 32'b0_000000_11110_00001_101_0100_0_1100011;  // bge x1, x30, 8

        //rom[x]=32'b imm20      _ rs1 _f3 _ rd  _ op // LU-Type, AU-Type
        rom[37] = 32'b00000000000000000001_00100_0110111;  // lui x4, 0x10000
        rom[38] = 32'b00000000000000000001_00101_0010111;  // auipc x5, 0x10000

        //rom[x]=32'b imm[20]_imm[10:1]_imm[11]_imm[19:12]_rd_op // J-Type
        rom[39] = 32'b0_0000000100_0_00000000_00110_1101111; // jal x6  PC 8증가.
        rom[40] = 32'b0000000_00000_00000_000_00000_0000000;

        //rom[x]=32'b imm12       _ rs1 _000 _ rd _  op // JL-Type, 
        rom[41] = 32'b000000000001_00001_000_00111_1100111; // jalr x7, x1, 1 PC 12증가.
        rom[42] = 32'b0000000_00000_00000_000_00000_0000000;
        rom[43] = 32'b0000000_00000_00000_000_00000_0000000;
        // 테스트용 R-Type add값 넣음.
        rom[44] = 32'b0000000_00001_00010_000_00111_0110011;
        */
    end

    assign data = rom[addr[31:2]];
endmodule

module twf1_2_rom (
  input  logic [8:0] addr,
  output logic signed [8:0] re,
  output logic signed [8:0] im
);

  wire signed [8:0] rom_re [0:511];
  wire signed [8:0] rom_im [0:511];

      assign rom_re[  0] =  128;    assign rom_im[  0] =    0;
      assign rom_re[  1] =  128;    assign rom_im[  1] =    0;
      assign rom_re[  2] =  128;    assign rom_im[  2] =    0;
      assign rom_re[  3] =  128;    assign rom_im[  3] =    0;
      assign rom_re[  4] =  128;    assign rom_im[  4] =    0;
      assign rom_re[  5] =  128;    assign rom_im[  5] =    0;
      assign rom_re[  6] =  128;    assign rom_im[  6] =    0;
      assign rom_re[  7] =  128;    assign rom_im[  7] =    0;
      assign rom_re[  8] =  128;    assign rom_im[  8] =    0;
      assign rom_re[  9] =  118;    assign rom_im[  9] =  -49;
      assign rom_re[ 10] =   91;    assign rom_im[ 10] =  -91;
      assign rom_re[ 11] =   49;    assign rom_im[ 11] = -118;
      assign rom_re[ 12] =    0;    assign rom_im[ 12] = -128;
      assign rom_re[ 13] =  -49;    assign rom_im[ 13] = -118;
      assign rom_re[ 14] =  -91;    assign rom_im[ 14] =  -91;
      assign rom_re[ 15] = -118;    assign rom_im[ 15] =  -49;
      assign rom_re[ 16] =  128;    assign rom_im[ 16] =    0;
      assign rom_re[ 17] =  126;    assign rom_im[ 17] =  -25;
      assign rom_re[ 18] =  118;    assign rom_im[ 18] =  -49;
      assign rom_re[ 19] =  106;    assign rom_im[ 19] =  -71;
      assign rom_re[ 20] =   91;    assign rom_im[ 20] =  -91;
      assign rom_re[ 21] =   71;    assign rom_im[ 21] = -106;
      assign rom_re[ 22] =   49;    assign rom_im[ 22] = -118;
      assign rom_re[ 23] =   25;    assign rom_im[ 23] = -126;
      assign rom_re[ 24] =  128;    assign rom_im[ 24] =    0;
      assign rom_re[ 25] =  106;    assign rom_im[ 25] =  -71;
      assign rom_re[ 26] =   49;    assign rom_im[ 26] = -118;
      assign rom_re[ 27] =  -25;    assign rom_im[ 27] = -126;
      assign rom_re[ 28] =  -91;    assign rom_im[ 28] =  -91;
      assign rom_re[ 29] = -126;    assign rom_im[ 29] =  -25;
      assign rom_re[ 30] = -118;    assign rom_im[ 30] =   49;
      assign rom_re[ 31] =  -71;    assign rom_im[ 31] =  106;
      assign rom_re[ 32] =  128;    assign rom_im[ 32] =    0;
      assign rom_re[ 33] =  127;    assign rom_im[ 33] =  -13;
      assign rom_re[ 34] =  126;    assign rom_im[ 34] =  -25;
      assign rom_re[ 35] =  122;    assign rom_im[ 35] =  -37;
      assign rom_re[ 36] =  118;    assign rom_im[ 36] =  -49;
      assign rom_re[ 37] =  113;    assign rom_im[ 37] =  -60;
      assign rom_re[ 38] =  106;    assign rom_im[ 38] =  -71;
      assign rom_re[ 39] =   99;    assign rom_im[ 39] =  -81;
      assign rom_re[ 40] =  128;    assign rom_im[ 40] =    0;
      assign rom_re[ 41] =  113;    assign rom_im[ 41] =  -60;
      assign rom_re[ 42] =   71;    assign rom_im[ 42] = -106;
      assign rom_re[ 43] =   13;    assign rom_im[ 43] = -127;
      assign rom_re[ 44] =  -49;    assign rom_im[ 44] = -118;
      assign rom_re[ 45] =  -99;    assign rom_im[ 45] =  -81;
      assign rom_re[ 46] = -126;    assign rom_im[ 46] =  -25;
      assign rom_re[ 47] = -122;    assign rom_im[ 47] =   37;
      assign rom_re[ 48] =  128;    assign rom_im[ 48] =    0;
      assign rom_re[ 49] =  122;    assign rom_im[ 49] =  -37;
      assign rom_re[ 50] =  106;    assign rom_im[ 50] =  -71;
      assign rom_re[ 51] =   81;    assign rom_im[ 51] =  -99;
      assign rom_re[ 52] =   49;    assign rom_im[ 52] = -118;
      assign rom_re[ 53] =   13;    assign rom_im[ 53] = -127;
      assign rom_re[ 54] =  -25;    assign rom_im[ 54] = -126;
      assign rom_re[ 55] =  -60;    assign rom_im[ 55] = -113;
      assign rom_re[ 56] =  128;    assign rom_im[ 56] =    0;
      assign rom_re[ 57] =   99;    assign rom_im[ 57] =  -81;
      assign rom_re[ 58] =   25;    assign rom_im[ 58] = -126;
      assign rom_re[ 59] =  -60;    assign rom_im[ 59] = -113;
      assign rom_re[ 60] = -118;    assign rom_im[ 60] =  -49;
      assign rom_re[ 61] = -122;    assign rom_im[ 61] =   37;
      assign rom_re[ 62] =  -71;    assign rom_im[ 62] =  106;
      assign rom_re[ 63] =   13;    assign rom_im[ 63] =  127;
      assign rom_re[ 64] =  128;    assign rom_im[ 64] =    0;
      assign rom_re[ 65] =  128;    assign rom_im[ 65] =    0;
      assign rom_re[ 66] =  128;    assign rom_im[ 66] =    0;
      assign rom_re[ 67] =  128;    assign rom_im[ 67] =    0;
      assign rom_re[ 68] =  128;    assign rom_im[ 68] =    0;
      assign rom_re[ 69] =  128;    assign rom_im[ 69] =    0;
      assign rom_re[ 70] =  128;    assign rom_im[ 70] =    0;
      assign rom_re[ 71] =  128;    assign rom_im[ 71] =    0;
      assign rom_re[ 72] =  128;    assign rom_im[ 72] =    0;
      assign rom_re[ 73] =  118;    assign rom_im[ 73] =  -49;
      assign rom_re[ 74] =   91;    assign rom_im[ 74] =  -91;
      assign rom_re[ 75] =   49;    assign rom_im[ 75] = -118;
      assign rom_re[ 76] =    0;    assign rom_im[ 76] = -128;
      assign rom_re[ 77] =  -49;    assign rom_im[ 77] = -118;
      assign rom_re[ 78] =  -91;    assign rom_im[ 78] =  -91;
      assign rom_re[ 79] = -118;    assign rom_im[ 79] =  -49;
      assign rom_re[ 80] =  128;    assign rom_im[ 80] =    0;
      assign rom_re[ 81] =  126;    assign rom_im[ 81] =  -25;
      assign rom_re[ 82] =  118;    assign rom_im[ 82] =  -49;
      assign rom_re[ 83] =  106;    assign rom_im[ 83] =  -71;
      assign rom_re[ 84] =   91;    assign rom_im[ 84] =  -91;
      assign rom_re[ 85] =   71;    assign rom_im[ 85] = -106;
      assign rom_re[ 86] =   49;    assign rom_im[ 86] = -118;
      assign rom_re[ 87] =   25;    assign rom_im[ 87] = -126;
      assign rom_re[ 88] =  128;    assign rom_im[ 88] =    0;
      assign rom_re[ 89] =  106;    assign rom_im[ 89] =  -71;
      assign rom_re[ 90] =   49;    assign rom_im[ 90] = -118;
      assign rom_re[ 91] =  -25;    assign rom_im[ 91] = -126;
      assign rom_re[ 92] =  -91;    assign rom_im[ 92] =  -91;
      assign rom_re[ 93] = -126;    assign rom_im[ 93] =  -25;
      assign rom_re[ 94] = -118;    assign rom_im[ 94] =   49;
      assign rom_re[ 95] =  -71;    assign rom_im[ 95] =  106;
      assign rom_re[ 96] =  128;    assign rom_im[ 96] =    0;
      assign rom_re[ 97] =  127;    assign rom_im[ 97] =  -13;
      assign rom_re[ 98] =  126;    assign rom_im[ 98] =  -25;
      assign rom_re[ 99] =  122;    assign rom_im[ 99] =  -37;
      assign rom_re[100] =  118;    assign rom_im[100] =  -49;
      assign rom_re[101] =  113;    assign rom_im[101] =  -60;
      assign rom_re[102] =  106;    assign rom_im[102] =  -71;
      assign rom_re[103] =   99;    assign rom_im[103] =  -81;
      assign rom_re[104] =  128;    assign rom_im[104] =    0;
      assign rom_re[105] =  113;    assign rom_im[105] =  -60;
      assign rom_re[106] =   71;    assign rom_im[106] = -106;
      assign rom_re[107] =   13;    assign rom_im[107] = -127;
      assign rom_re[108] =  -49;    assign rom_im[108] = -118;
      assign rom_re[109] =  -99;    assign rom_im[109] =  -81;
      assign rom_re[110] = -126;    assign rom_im[110] =  -25;
      assign rom_re[111] = -122;    assign rom_im[111] =   37;
      assign rom_re[112] =  128;    assign rom_im[112] =    0;
      assign rom_re[113] =  122;    assign rom_im[113] =  -37;
      assign rom_re[114] =  106;    assign rom_im[114] =  -71;
      assign rom_re[115] =   81;    assign rom_im[115] =  -99;
      assign rom_re[116] =   49;    assign rom_im[116] = -118;
      assign rom_re[117] =   13;    assign rom_im[117] = -127;
      assign rom_re[118] =  -25;    assign rom_im[118] = -126;
      assign rom_re[119] =  -60;    assign rom_im[119] = -113;
      assign rom_re[120] =  128;    assign rom_im[120] =    0;
      assign rom_re[121] =   99;    assign rom_im[121] =  -81;
      assign rom_re[122] =   25;    assign rom_im[122] = -126;
      assign rom_re[123] =  -60;    assign rom_im[123] = -113;
      assign rom_re[124] = -118;    assign rom_im[124] =  -49;
      assign rom_re[125] = -122;    assign rom_im[125] =   37;
      assign rom_re[126] =  -71;    assign rom_im[126] =  106;
      assign rom_re[127] =   13;    assign rom_im[127] =  127;
      assign rom_re[128] =  128;    assign rom_im[128] =    0;
      assign rom_re[129] =  128;    assign rom_im[129] =    0;
      assign rom_re[130] =  128;    assign rom_im[130] =    0;
      assign rom_re[131] =  128;    assign rom_im[131] =    0;
      assign rom_re[132] =  128;    assign rom_im[132] =    0;
      assign rom_re[133] =  128;    assign rom_im[133] =    0;
      assign rom_re[134] =  128;    assign rom_im[134] =    0;
      assign rom_re[135] =  128;    assign rom_im[135] =    0;
      assign rom_re[136] =  128;    assign rom_im[136] =    0;
      assign rom_re[137] =  118;    assign rom_im[137] =  -49;
      assign rom_re[138] =   91;    assign rom_im[138] =  -91;
      assign rom_re[139] =   49;    assign rom_im[139] = -118;
      assign rom_re[140] =    0;    assign rom_im[140] = -128;
      assign rom_re[141] =  -49;    assign rom_im[141] = -118;
      assign rom_re[142] =  -91;    assign rom_im[142] =  -91;
      assign rom_re[143] = -118;    assign rom_im[143] =  -49;
      assign rom_re[144] =  128;    assign rom_im[144] =    0;
      assign rom_re[145] =  126;    assign rom_im[145] =  -25;
      assign rom_re[146] =  118;    assign rom_im[146] =  -49;
      assign rom_re[147] =  106;    assign rom_im[147] =  -71;
      assign rom_re[148] =   91;    assign rom_im[148] =  -91;
      assign rom_re[149] =   71;    assign rom_im[149] = -106;
      assign rom_re[150] =   49;    assign rom_im[150] = -118;
      assign rom_re[151] =   25;    assign rom_im[151] = -126;
      assign rom_re[152] =  128;    assign rom_im[152] =    0;
      assign rom_re[153] =  106;    assign rom_im[153] =  -71;
      assign rom_re[154] =   49;    assign rom_im[154] = -118;
      assign rom_re[155] =  -25;    assign rom_im[155] = -126;
      assign rom_re[156] =  -91;    assign rom_im[156] =  -91;
      assign rom_re[157] = -126;    assign rom_im[157] =  -25;
      assign rom_re[158] = -118;    assign rom_im[158] =   49;
      assign rom_re[159] =  -71;    assign rom_im[159] =  106;
      assign rom_re[160] =  128;    assign rom_im[160] =    0;
      assign rom_re[161] =  127;    assign rom_im[161] =  -13;
      assign rom_re[162] =  126;    assign rom_im[162] =  -25;
      assign rom_re[163] =  122;    assign rom_im[163] =  -37;
      assign rom_re[164] =  118;    assign rom_im[164] =  -49;
      assign rom_re[165] =  113;    assign rom_im[165] =  -60;
      assign rom_re[166] =  106;    assign rom_im[166] =  -71;
      assign rom_re[167] =   99;    assign rom_im[167] =  -81;
      assign rom_re[168] =  128;    assign rom_im[168] =    0;
      assign rom_re[169] =  113;    assign rom_im[169] =  -60;
      assign rom_re[170] =   71;    assign rom_im[170] = -106;
      assign rom_re[171] =   13;    assign rom_im[171] = -127;
      assign rom_re[172] =  -49;    assign rom_im[172] = -118;
      assign rom_re[173] =  -99;    assign rom_im[173] =  -81;
      assign rom_re[174] = -126;    assign rom_im[174] =  -25;
      assign rom_re[175] = -122;    assign rom_im[175] =   37;
      assign rom_re[176] =  128;    assign rom_im[176] =    0;
      assign rom_re[177] =  122;    assign rom_im[177] =  -37;
      assign rom_re[178] =  106;    assign rom_im[178] =  -71;
      assign rom_re[179] =   81;    assign rom_im[179] =  -99;
      assign rom_re[180] =   49;    assign rom_im[180] = -118;
      assign rom_re[181] =   13;    assign rom_im[181] = -127;
      assign rom_re[182] =  -25;    assign rom_im[182] = -126;
      assign rom_re[183] =  -60;    assign rom_im[183] = -113;
      assign rom_re[184] =  128;    assign rom_im[184] =    0;
      assign rom_re[185] =   99;    assign rom_im[185] =  -81;
      assign rom_re[186] =   25;    assign rom_im[186] = -126;
      assign rom_re[187] =  -60;    assign rom_im[187] = -113;
      assign rom_re[188] = -118;    assign rom_im[188] =  -49;
      assign rom_re[189] = -122;    assign rom_im[189] =   37;
      assign rom_re[190] =  -71;    assign rom_im[190] =  106;
      assign rom_re[191] =   13;    assign rom_im[191] =  127;
      assign rom_re[192] =  128;    assign rom_im[192] =    0;
      assign rom_re[193] =  128;    assign rom_im[193] =    0;
      assign rom_re[194] =  128;    assign rom_im[194] =    0;
      assign rom_re[195] =  128;    assign rom_im[195] =    0;
      assign rom_re[196] =  128;    assign rom_im[196] =    0;
      assign rom_re[197] =  128;    assign rom_im[197] =    0;
      assign rom_re[198] =  128;    assign rom_im[198] =    0;
      assign rom_re[199] =  128;    assign rom_im[199] =    0;
      assign rom_re[200] =  128;    assign rom_im[200] =    0;
      assign rom_re[201] =  118;    assign rom_im[201] =  -49;
      assign rom_re[202] =   91;    assign rom_im[202] =  -91;
      assign rom_re[203] =   49;    assign rom_im[203] = -118;
      assign rom_re[204] =    0;    assign rom_im[204] = -128;
      assign rom_re[205] =  -49;    assign rom_im[205] = -118;
      assign rom_re[206] =  -91;    assign rom_im[206] =  -91;
      assign rom_re[207] = -118;    assign rom_im[207] =  -49;
      assign rom_re[208] =  128;    assign rom_im[208] =    0;
      assign rom_re[209] =  126;    assign rom_im[209] =  -25;
      assign rom_re[210] =  118;    assign rom_im[210] =  -49;
      assign rom_re[211] =  106;    assign rom_im[211] =  -71;
      assign rom_re[212] =   91;    assign rom_im[212] =  -91;
      assign rom_re[213] =   71;    assign rom_im[213] = -106;
      assign rom_re[214] =   49;    assign rom_im[214] = -118;
      assign rom_re[215] =   25;    assign rom_im[215] = -126;
      assign rom_re[216] =  128;    assign rom_im[216] =    0;
      assign rom_re[217] =  106;    assign rom_im[217] =  -71;
      assign rom_re[218] =   49;    assign rom_im[218] = -118;
      assign rom_re[219] =  -25;    assign rom_im[219] = -126;
      assign rom_re[220] =  -91;    assign rom_im[220] =  -91;
      assign rom_re[221] = -126;    assign rom_im[221] =  -25;
      assign rom_re[222] = -118;    assign rom_im[222] =   49;
      assign rom_re[223] =  -71;    assign rom_im[223] =  106;
      assign rom_re[224] =  128;    assign rom_im[224] =    0;
      assign rom_re[225] =  127;    assign rom_im[225] =  -13;
      assign rom_re[226] =  126;    assign rom_im[226] =  -25;
      assign rom_re[227] =  122;    assign rom_im[227] =  -37;
      assign rom_re[228] =  118;    assign rom_im[228] =  -49;
      assign rom_re[229] =  113;    assign rom_im[229] =  -60;
      assign rom_re[230] =  106;    assign rom_im[230] =  -71;
      assign rom_re[231] =   99;    assign rom_im[231] =  -81;
      assign rom_re[232] =  128;    assign rom_im[232] =    0;
      assign rom_re[233] =  113;    assign rom_im[233] =  -60;
      assign rom_re[234] =   71;    assign rom_im[234] = -106;
      assign rom_re[235] =   13;    assign rom_im[235] = -127;
      assign rom_re[236] =  -49;    assign rom_im[236] = -118;
      assign rom_re[237] =  -99;    assign rom_im[237] =  -81;
      assign rom_re[238] = -126;    assign rom_im[238] =  -25;
      assign rom_re[239] = -122;    assign rom_im[239] =   37;
      assign rom_re[240] =  128;    assign rom_im[240] =    0;
      assign rom_re[241] =  122;    assign rom_im[241] =  -37;
      assign rom_re[242] =  106;    assign rom_im[242] =  -71;
      assign rom_re[243] =   81;    assign rom_im[243] =  -99;
      assign rom_re[244] =   49;    assign rom_im[244] = -118;
      assign rom_re[245] =   13;    assign rom_im[245] = -127;
      assign rom_re[246] =  -25;    assign rom_im[246] = -126;
      assign rom_re[247] =  -60;    assign rom_im[247] = -113;
      assign rom_re[248] =  128;    assign rom_im[248] =    0;
      assign rom_re[249] =   99;    assign rom_im[249] =  -81;
      assign rom_re[250] =   25;    assign rom_im[250] = -126;
      assign rom_re[251] =  -60;    assign rom_im[251] = -113;
      assign rom_re[252] = -118;    assign rom_im[252] =  -49;
      assign rom_re[253] = -122;    assign rom_im[253] =   37;
      assign rom_re[254] =  -71;    assign rom_im[254] =  106;
      assign rom_re[255] =   13;    assign rom_im[255] =  127;
      assign rom_re[256] =  128;    assign rom_im[256] =    0;
      assign rom_re[257] =  128;    assign rom_im[257] =    0;
      assign rom_re[258] =  128;    assign rom_im[258] =    0;
      assign rom_re[259] =  128;    assign rom_im[259] =    0;
      assign rom_re[260] =  128;    assign rom_im[260] =    0;
      assign rom_re[261] =  128;    assign rom_im[261] =    0;
      assign rom_re[262] =  128;    assign rom_im[262] =    0;
      assign rom_re[263] =  128;    assign rom_im[263] =    0;
      assign rom_re[264] =  128;    assign rom_im[264] =    0;
      assign rom_re[265] =  118;    assign rom_im[265] =  -49;
      assign rom_re[266] =   91;    assign rom_im[266] =  -91;
      assign rom_re[267] =   49;    assign rom_im[267] = -118;
      assign rom_re[268] =    0;    assign rom_im[268] = -128;
      assign rom_re[269] =  -49;    assign rom_im[269] = -118;
      assign rom_re[270] =  -91;    assign rom_im[270] =  -91;
      assign rom_re[271] = -118;    assign rom_im[271] =  -49;
      assign rom_re[272] =  128;    assign rom_im[272] =    0;
      assign rom_re[273] =  126;    assign rom_im[273] =  -25;
      assign rom_re[274] =  118;    assign rom_im[274] =  -49;
      assign rom_re[275] =  106;    assign rom_im[275] =  -71;
      assign rom_re[276] =   91;    assign rom_im[276] =  -91;
      assign rom_re[277] =   71;    assign rom_im[277] = -106;
      assign rom_re[278] =   49;    assign rom_im[278] = -118;
      assign rom_re[279] =   25;    assign rom_im[279] = -126;
      assign rom_re[280] =  128;    assign rom_im[280] =    0;
      assign rom_re[281] =  106;    assign rom_im[281] =  -71;
      assign rom_re[282] =   49;    assign rom_im[282] = -118;
      assign rom_re[283] =  -25;    assign rom_im[283] = -126;
      assign rom_re[284] =  -91;    assign rom_im[284] =  -91;
      assign rom_re[285] = -126;    assign rom_im[285] =  -25;
      assign rom_re[286] = -118;    assign rom_im[286] =   49;
      assign rom_re[287] =  -71;    assign rom_im[287] =  106;
      assign rom_re[288] =  128;    assign rom_im[288] =    0;
      assign rom_re[289] =  127;    assign rom_im[289] =  -13;
      assign rom_re[290] =  126;    assign rom_im[290] =  -25;
      assign rom_re[291] =  122;    assign rom_im[291] =  -37;
      assign rom_re[292] =  118;    assign rom_im[292] =  -49;
      assign rom_re[293] =  113;    assign rom_im[293] =  -60;
      assign rom_re[294] =  106;    assign rom_im[294] =  -71;
      assign rom_re[295] =   99;    assign rom_im[295] =  -81;
      assign rom_re[296] =  128;    assign rom_im[296] =    0;
      assign rom_re[297] =  113;    assign rom_im[297] =  -60;
      assign rom_re[298] =   71;    assign rom_im[298] = -106;
      assign rom_re[299] =   13;    assign rom_im[299] = -127;
      assign rom_re[300] =  -49;    assign rom_im[300] = -118;
      assign rom_re[301] =  -99;    assign rom_im[301] =  -81;
      assign rom_re[302] = -126;    assign rom_im[302] =  -25;
      assign rom_re[303] = -122;    assign rom_im[303] =   37;
      assign rom_re[304] =  128;    assign rom_im[304] =    0;
      assign rom_re[305] =  122;    assign rom_im[305] =  -37;
      assign rom_re[306] =  106;    assign rom_im[306] =  -71;
      assign rom_re[307] =   81;    assign rom_im[307] =  -99;
      assign rom_re[308] =   49;    assign rom_im[308] = -118;
      assign rom_re[309] =   13;    assign rom_im[309] = -127;
      assign rom_re[310] =  -25;    assign rom_im[310] = -126;
      assign rom_re[311] =  -60;    assign rom_im[311] = -113;
      assign rom_re[312] =  128;    assign rom_im[312] =    0;
      assign rom_re[313] =   99;    assign rom_im[313] =  -81;
      assign rom_re[314] =   25;    assign rom_im[314] = -126;
      assign rom_re[315] =  -60;    assign rom_im[315] = -113;
      assign rom_re[316] = -118;    assign rom_im[316] =  -49;
      assign rom_re[317] = -122;    assign rom_im[317] =   37;
      assign rom_re[318] =  -71;    assign rom_im[318] =  106;
      assign rom_re[319] =   13;    assign rom_im[319] =  127;
      assign rom_re[320] =  128;    assign rom_im[320] =    0;
      assign rom_re[321] =  128;    assign rom_im[321] =    0;
      assign rom_re[322] =  128;    assign rom_im[322] =    0;
      assign rom_re[323] =  128;    assign rom_im[323] =    0;
      assign rom_re[324] =  128;    assign rom_im[324] =    0;
      assign rom_re[325] =  128;    assign rom_im[325] =    0;
      assign rom_re[326] =  128;    assign rom_im[326] =    0;
      assign rom_re[327] =  128;    assign rom_im[327] =    0;
      assign rom_re[328] =  128;    assign rom_im[328] =    0;
      assign rom_re[329] =  118;    assign rom_im[329] =  -49;
      assign rom_re[330] =   91;    assign rom_im[330] =  -91;
      assign rom_re[331] =   49;    assign rom_im[331] = -118;
      assign rom_re[332] =    0;    assign rom_im[332] = -128;
      assign rom_re[333] =  -49;    assign rom_im[333] = -118;
      assign rom_re[334] =  -91;    assign rom_im[334] =  -91;
      assign rom_re[335] = -118;    assign rom_im[335] =  -49;
      assign rom_re[336] =  128;    assign rom_im[336] =    0;
      assign rom_re[337] =  126;    assign rom_im[337] =  -25;
      assign rom_re[338] =  118;    assign rom_im[338] =  -49;
      assign rom_re[339] =  106;    assign rom_im[339] =  -71;
      assign rom_re[340] =   91;    assign rom_im[340] =  -91;
      assign rom_re[341] =   71;    assign rom_im[341] = -106;
      assign rom_re[342] =   49;    assign rom_im[342] = -118;
      assign rom_re[343] =   25;    assign rom_im[343] = -126;
      assign rom_re[344] =  128;    assign rom_im[344] =    0;
      assign rom_re[345] =  106;    assign rom_im[345] =  -71;
      assign rom_re[346] =   49;    assign rom_im[346] = -118;
      assign rom_re[347] =  -25;    assign rom_im[347] = -126;
      assign rom_re[348] =  -91;    assign rom_im[348] =  -91;
      assign rom_re[349] = -126;    assign rom_im[349] =  -25;
      assign rom_re[350] = -118;    assign rom_im[350] =   49;
      assign rom_re[351] =  -71;    assign rom_im[351] =  106;
      assign rom_re[352] =  128;    assign rom_im[352] =    0;
      assign rom_re[353] =  127;    assign rom_im[353] =  -13;
      assign rom_re[354] =  126;    assign rom_im[354] =  -25;
      assign rom_re[355] =  122;    assign rom_im[355] =  -37;
      assign rom_re[356] =  118;    assign rom_im[356] =  -49;
      assign rom_re[357] =  113;    assign rom_im[357] =  -60;
      assign rom_re[358] =  106;    assign rom_im[358] =  -71;
      assign rom_re[359] =   99;    assign rom_im[359] =  -81;
      assign rom_re[360] =  128;    assign rom_im[360] =    0;
      assign rom_re[361] =  113;    assign rom_im[361] =  -60;
      assign rom_re[362] =   71;    assign rom_im[362] = -106;
      assign rom_re[363] =   13;    assign rom_im[363] = -127;
      assign rom_re[364] =  -49;    assign rom_im[364] = -118;
      assign rom_re[365] =  -99;    assign rom_im[365] =  -81;
      assign rom_re[366] = -126;    assign rom_im[366] =  -25;
      assign rom_re[367] = -122;    assign rom_im[367] =   37;
      assign rom_re[368] =  128;    assign rom_im[368] =    0;
      assign rom_re[369] =  122;    assign rom_im[369] =  -37;
      assign rom_re[370] =  106;    assign rom_im[370] =  -71;
      assign rom_re[371] =   81;    assign rom_im[371] =  -99;
      assign rom_re[372] =   49;    assign rom_im[372] = -118;
      assign rom_re[373] =   13;    assign rom_im[373] = -127;
      assign rom_re[374] =  -25;    assign rom_im[374] = -126;
      assign rom_re[375] =  -60;    assign rom_im[375] = -113;
      assign rom_re[376] =  128;    assign rom_im[376] =    0;
      assign rom_re[377] =   99;    assign rom_im[377] =  -81;
      assign rom_re[378] =   25;    assign rom_im[378] = -126;
      assign rom_re[379] =  -60;    assign rom_im[379] = -113;
      assign rom_re[380] = -118;    assign rom_im[380] =  -49;
      assign rom_re[381] = -122;    assign rom_im[381] =   37;
      assign rom_re[382] =  -71;    assign rom_im[382] =  106;
      assign rom_re[383] =   13;    assign rom_im[383] =  127;
      assign rom_re[384] =  128;    assign rom_im[384] =    0;
      assign rom_re[385] =  128;    assign rom_im[385] =    0;
      assign rom_re[386] =  128;    assign rom_im[386] =    0;
      assign rom_re[387] =  128;    assign rom_im[387] =    0;
      assign rom_re[388] =  128;    assign rom_im[388] =    0;
      assign rom_re[389] =  128;    assign rom_im[389] =    0;
      assign rom_re[390] =  128;    assign rom_im[390] =    0;
      assign rom_re[391] =  128;    assign rom_im[391] =    0;
      assign rom_re[392] =  128;    assign rom_im[392] =    0;
      assign rom_re[393] =  118;    assign rom_im[393] =  -49;
      assign rom_re[394] =   91;    assign rom_im[394] =  -91;
      assign rom_re[395] =   49;    assign rom_im[395] = -118;
      assign rom_re[396] =    0;    assign rom_im[396] = -128;
      assign rom_re[397] =  -49;    assign rom_im[397] = -118;
      assign rom_re[398] =  -91;    assign rom_im[398] =  -91;
      assign rom_re[399] = -118;    assign rom_im[399] =  -49;
      assign rom_re[400] =  128;    assign rom_im[400] =    0;
      assign rom_re[401] =  126;    assign rom_im[401] =  -25;
      assign rom_re[402] =  118;    assign rom_im[402] =  -49;
      assign rom_re[403] =  106;    assign rom_im[403] =  -71;
      assign rom_re[404] =   91;    assign rom_im[404] =  -91;
      assign rom_re[405] =   71;    assign rom_im[405] = -106;
      assign rom_re[406] =   49;    assign rom_im[406] = -118;
      assign rom_re[407] =   25;    assign rom_im[407] = -126;
      assign rom_re[408] =  128;    assign rom_im[408] =    0;
      assign rom_re[409] =  106;    assign rom_im[409] =  -71;
      assign rom_re[410] =   49;    assign rom_im[410] = -118;
      assign rom_re[411] =  -25;    assign rom_im[411] = -126;
      assign rom_re[412] =  -91;    assign rom_im[412] =  -91;
      assign rom_re[413] = -126;    assign rom_im[413] =  -25;
      assign rom_re[414] = -118;    assign rom_im[414] =   49;
      assign rom_re[415] =  -71;    assign rom_im[415] =  106;
      assign rom_re[416] =  128;    assign rom_im[416] =    0;
      assign rom_re[417] =  127;    assign rom_im[417] =  -13;
      assign rom_re[418] =  126;    assign rom_im[418] =  -25;
      assign rom_re[419] =  122;    assign rom_im[419] =  -37;
      assign rom_re[420] =  118;    assign rom_im[420] =  -49;
      assign rom_re[421] =  113;    assign rom_im[421] =  -60;
      assign rom_re[422] =  106;    assign rom_im[422] =  -71;
      assign rom_re[423] =   99;    assign rom_im[423] =  -81;
      assign rom_re[424] =  128;    assign rom_im[424] =    0;
      assign rom_re[425] =  113;    assign rom_im[425] =  -60;
      assign rom_re[426] =   71;    assign rom_im[426] = -106;
      assign rom_re[427] =   13;    assign rom_im[427] = -127;
      assign rom_re[428] =  -49;    assign rom_im[428] = -118;
      assign rom_re[429] =  -99;    assign rom_im[429] =  -81;
      assign rom_re[430] = -126;    assign rom_im[430] =  -25;
      assign rom_re[431] = -122;    assign rom_im[431] =   37;
      assign rom_re[432] =  128;    assign rom_im[432] =    0;
      assign rom_re[433] =  122;    assign rom_im[433] =  -37;
      assign rom_re[434] =  106;    assign rom_im[434] =  -71;
      assign rom_re[435] =   81;    assign rom_im[435] =  -99;
      assign rom_re[436] =   49;    assign rom_im[436] = -118;
      assign rom_re[437] =   13;    assign rom_im[437] = -127;
      assign rom_re[438] =  -25;    assign rom_im[438] = -126;
      assign rom_re[439] =  -60;    assign rom_im[439] = -113;
      assign rom_re[440] =  128;    assign rom_im[440] =    0;
      assign rom_re[441] =   99;    assign rom_im[441] =  -81;
      assign rom_re[442] =   25;    assign rom_im[442] = -126;
      assign rom_re[443] =  -60;    assign rom_im[443] = -113;
      assign rom_re[444] = -118;    assign rom_im[444] =  -49;
      assign rom_re[445] = -122;    assign rom_im[445] =   37;
      assign rom_re[446] =  -71;    assign rom_im[446] =  106;
      assign rom_re[447] =   13;    assign rom_im[447] =  127;
      assign rom_re[448] =  128;    assign rom_im[448] =    0;
      assign rom_re[449] =  128;    assign rom_im[449] =    0;
      assign rom_re[450] =  128;    assign rom_im[450] =    0;
      assign rom_re[451] =  128;    assign rom_im[451] =    0;
      assign rom_re[452] =  128;    assign rom_im[452] =    0;
      assign rom_re[453] =  128;    assign rom_im[453] =    0;
      assign rom_re[454] =  128;    assign rom_im[454] =    0;
      assign rom_re[455] =  128;    assign rom_im[455] =    0;
      assign rom_re[456] =  128;    assign rom_im[456] =    0;
      assign rom_re[457] =  118;    assign rom_im[457] =  -49;
      assign rom_re[458] =   91;    assign rom_im[458] =  -91;
      assign rom_re[459] =   49;    assign rom_im[459] = -118;
      assign rom_re[460] =    0;    assign rom_im[460] = -128;
      assign rom_re[461] =  -49;    assign rom_im[461] = -118;
      assign rom_re[462] =  -91;    assign rom_im[462] =  -91;
      assign rom_re[463] = -118;    assign rom_im[463] =  -49;
      assign rom_re[464] =  128;    assign rom_im[464] =    0;
      assign rom_re[465] =  126;    assign rom_im[465] =  -25;
      assign rom_re[466] =  118;    assign rom_im[466] =  -49;
      assign rom_re[467] =  106;    assign rom_im[467] =  -71;
      assign rom_re[468] =   91;    assign rom_im[468] =  -91;
      assign rom_re[469] =   71;    assign rom_im[469] = -106;
      assign rom_re[470] =   49;    assign rom_im[470] = -118;
      assign rom_re[471] =   25;    assign rom_im[471] = -126;
      assign rom_re[472] =  128;    assign rom_im[472] =    0;
      assign rom_re[473] =  106;    assign rom_im[473] =  -71;
      assign rom_re[474] =   49;    assign rom_im[474] = -118;
      assign rom_re[475] =  -25;    assign rom_im[475] = -126;
      assign rom_re[476] =  -91;    assign rom_im[476] =  -91;
      assign rom_re[477] = -126;    assign rom_im[477] =  -25;
      assign rom_re[478] = -118;    assign rom_im[478] =   49;
      assign rom_re[479] =  -71;    assign rom_im[479] =  106;
      assign rom_re[480] =  128;    assign rom_im[480] =    0;
      assign rom_re[481] =  127;    assign rom_im[481] =  -13;
      assign rom_re[482] =  126;    assign rom_im[482] =  -25;
      assign rom_re[483] =  122;    assign rom_im[483] =  -37;
      assign rom_re[484] =  118;    assign rom_im[484] =  -49;
      assign rom_re[485] =  113;    assign rom_im[485] =  -60;
      assign rom_re[486] =  106;    assign rom_im[486] =  -71;
      assign rom_re[487] =   99;    assign rom_im[487] =  -81;
      assign rom_re[488] =  128;    assign rom_im[488] =    0;
      assign rom_re[489] =  113;    assign rom_im[489] =  -60;
      assign rom_re[490] =   71;    assign rom_im[490] = -106;
      assign rom_re[491] =   13;    assign rom_im[491] = -127;
      assign rom_re[492] =  -49;    assign rom_im[492] = -118;
      assign rom_re[493] =  -99;    assign rom_im[493] =  -81;
      assign rom_re[494] = -126;    assign rom_im[494] =  -25;
      assign rom_re[495] = -122;    assign rom_im[495] =   37;
      assign rom_re[496] =  128;    assign rom_im[496] =    0;
      assign rom_re[497] =  122;    assign rom_im[497] =  -37;
      assign rom_re[498] =  106;    assign rom_im[498] =  -71;
      assign rom_re[499] =   81;    assign rom_im[499] =  -99;
      assign rom_re[500] =   49;    assign rom_im[500] = -118;
      assign rom_re[501] =   13;    assign rom_im[501] = -127;
      assign rom_re[502] =  -25;    assign rom_im[502] = -126;
      assign rom_re[503] =  -60;    assign rom_im[503] = -113;
      assign rom_re[504] =  128;    assign rom_im[504] =    0;
      assign rom_re[505] =   99;    assign rom_im[505] =  -81;
      assign rom_re[506] =   25;    assign rom_im[506] = -126;
      assign rom_re[507] =  -60;    assign rom_im[507] = -113;
      assign rom_re[508] = -118;    assign rom_im[508] =  -49;
      assign rom_re[509] = -122;    assign rom_im[509] =   37;
      assign rom_re[510] =  -71;    assign rom_im[510] =  106;
      assign rom_re[511] =   13;    assign rom_im[511] =  127;

  assign re = rom_re[addr];
  assign im = rom_im[addr];

endmodule

module twf2_1_rom (
  input  logic [8:0] addr, // 0 ~ 511 address
  output logic signed [9:0] re,
  output logic signed [9:0] im
);

  wire signed [9:0] rom_re [511:0];
  wire signed [9:0] rom_im [511:0];
	
  assign re = rom_re[addr];
  assign im = rom_im[addr];

      assign rom_re[  0] =  256;    assign rom_im[  0] =    0;
      assign rom_re[  1] =  256;    assign rom_im[  1] =    0;
      assign rom_re[  2] =  256;    assign rom_im[  2] =    0;
      assign rom_re[  3] =    0;    assign rom_im[  3] = -256;
      assign rom_re[  4] =  256;    assign rom_im[  4] =    0;
      assign rom_re[  5] =  181;    assign rom_im[  5] = -181;
      assign rom_re[  6] =  256;    assign rom_im[  6] =    0;
      assign rom_re[  7] = -181;    assign rom_im[  7] = -181;
      assign rom_re[  8] =  256;    assign rom_im[  8] =    0;
      assign rom_re[  9] =  256;    assign rom_im[  9] =    0;
      assign rom_re[ 10] =  256;    assign rom_im[ 10] =    0;
      assign rom_re[ 11] =    0;    assign rom_im[ 11] = -256;
      assign rom_re[ 12] =  256;    assign rom_im[ 12] =    0;
      assign rom_re[ 13] =  181;    assign rom_im[ 13] = -181;
      assign rom_re[ 14] =  256;    assign rom_im[ 14] =    0;
      assign rom_re[ 15] = -181;    assign rom_im[ 15] = -181;
      assign rom_re[ 16] =  256;    assign rom_im[ 16] =    0;
      assign rom_re[ 17] =  256;    assign rom_im[ 17] =    0;
      assign rom_re[ 18] =  256;    assign rom_im[ 18] =    0;
      assign rom_re[ 19] =    0;    assign rom_im[ 19] = -256;
      assign rom_re[ 20] =  256;    assign rom_im[ 20] =    0;
      assign rom_re[ 21] =  181;    assign rom_im[ 21] = -181;
      assign rom_re[ 22] =  256;    assign rom_im[ 22] =    0;
      assign rom_re[ 23] = -181;    assign rom_im[ 23] = -181;
      assign rom_re[ 24] =  256;    assign rom_im[ 24] =    0;
      assign rom_re[ 25] =  256;    assign rom_im[ 25] =    0;
      assign rom_re[ 26] =  256;    assign rom_im[ 26] =    0;
      assign rom_re[ 27] =    0;    assign rom_im[ 27] = -256;
      assign rom_re[ 28] =  256;    assign rom_im[ 28] =    0;
      assign rom_re[ 29] =  181;    assign rom_im[ 29] = -181;
      assign rom_re[ 30] =  256;    assign rom_im[ 30] =    0;
      assign rom_re[ 31] = -181;    assign rom_im[ 31] = -181;
      assign rom_re[ 32] =  256;    assign rom_im[ 32] =    0;
      assign rom_re[ 33] =  256;    assign rom_im[ 33] =    0;
      assign rom_re[ 34] =  256;    assign rom_im[ 34] =    0;
      assign rom_re[ 35] =    0;    assign rom_im[ 35] = -256;
      assign rom_re[ 36] =  256;    assign rom_im[ 36] =    0;
      assign rom_re[ 37] =  181;    assign rom_im[ 37] = -181;
      assign rom_re[ 38] =  256;    assign rom_im[ 38] =    0;
      assign rom_re[ 39] = -181;    assign rom_im[ 39] = -181;
      assign rom_re[ 40] =  256;    assign rom_im[ 40] =    0;
      assign rom_re[ 41] =  256;    assign rom_im[ 41] =    0;
      assign rom_re[ 42] =  256;    assign rom_im[ 42] =    0;
      assign rom_re[ 43] =    0;    assign rom_im[ 43] = -256;
      assign rom_re[ 44] =  256;    assign rom_im[ 44] =    0;
      assign rom_re[ 45] =  181;    assign rom_im[ 45] = -181;
      assign rom_re[ 46] =  256;    assign rom_im[ 46] =    0;
      assign rom_re[ 47] = -181;    assign rom_im[ 47] = -181;
      assign rom_re[ 48] =  256;    assign rom_im[ 48] =    0;
      assign rom_re[ 49] =  256;    assign rom_im[ 49] =    0;
      assign rom_re[ 50] =  256;    assign rom_im[ 50] =    0;
      assign rom_re[ 51] =    0;    assign rom_im[ 51] = -256;
      assign rom_re[ 52] =  256;    assign rom_im[ 52] =    0;
      assign rom_re[ 53] =  181;    assign rom_im[ 53] = -181;
      assign rom_re[ 54] =  256;    assign rom_im[ 54] =    0;
      assign rom_re[ 55] = -181;    assign rom_im[ 55] = -181;
      assign rom_re[ 56] =  256;    assign rom_im[ 56] =    0;
      assign rom_re[ 57] =  256;    assign rom_im[ 57] =    0;
      assign rom_re[ 58] =  256;    assign rom_im[ 58] =    0;
      assign rom_re[ 59] =    0;    assign rom_im[ 59] = -256;
      assign rom_re[ 60] =  256;    assign rom_im[ 60] =    0;
      assign rom_re[ 61] =  181;    assign rom_im[ 61] = -181;
      assign rom_re[ 62] =  256;    assign rom_im[ 62] =    0;
      assign rom_re[ 63] = -181;    assign rom_im[ 63] = -181;
      assign rom_re[ 64] =  256;    assign rom_im[ 64] =    0;
      assign rom_re[ 65] =  256;    assign rom_im[ 65] =    0;
      assign rom_re[ 66] =  256;    assign rom_im[ 66] =    0;
      assign rom_re[ 67] =    0;    assign rom_im[ 67] = -256;
      assign rom_re[ 68] =  256;    assign rom_im[ 68] =    0;
      assign rom_re[ 69] =  181;    assign rom_im[ 69] = -181;
      assign rom_re[ 70] =  256;    assign rom_im[ 70] =    0;
      assign rom_re[ 71] = -181;    assign rom_im[ 71] = -181;
      assign rom_re[ 72] =  256;    assign rom_im[ 72] =    0;
      assign rom_re[ 73] =  256;    assign rom_im[ 73] =    0;
      assign rom_re[ 74] =  256;    assign rom_im[ 74] =    0;
      assign rom_re[ 75] =    0;    assign rom_im[ 75] = -256;
      assign rom_re[ 76] =  256;    assign rom_im[ 76] =    0;
      assign rom_re[ 77] =  181;    assign rom_im[ 77] = -181;
      assign rom_re[ 78] =  256;    assign rom_im[ 78] =    0;
      assign rom_re[ 79] = -181;    assign rom_im[ 79] = -181;
      assign rom_re[ 80] =  256;    assign rom_im[ 80] =    0;
      assign rom_re[ 81] =  256;    assign rom_im[ 81] =    0;
      assign rom_re[ 82] =  256;    assign rom_im[ 82] =    0;
      assign rom_re[ 83] =    0;    assign rom_im[ 83] = -256;
      assign rom_re[ 84] =  256;    assign rom_im[ 84] =    0;
      assign rom_re[ 85] =  181;    assign rom_im[ 85] = -181;
      assign rom_re[ 86] =  256;    assign rom_im[ 86] =    0;
      assign rom_re[ 87] = -181;    assign rom_im[ 87] = -181;
      assign rom_re[ 88] =  256;    assign rom_im[ 88] =    0;
      assign rom_re[ 89] =  256;    assign rom_im[ 89] =    0;
      assign rom_re[ 90] =  256;    assign rom_im[ 90] =    0;
      assign rom_re[ 91] =    0;    assign rom_im[ 91] = -256;
      assign rom_re[ 92] =  256;    assign rom_im[ 92] =    0;
      assign rom_re[ 93] =  181;    assign rom_im[ 93] = -181;
      assign rom_re[ 94] =  256;    assign rom_im[ 94] =    0;
      assign rom_re[ 95] = -181;    assign rom_im[ 95] = -181;
      assign rom_re[ 96] =  256;    assign rom_im[ 96] =    0;
      assign rom_re[ 97] =  256;    assign rom_im[ 97] =    0;
      assign rom_re[ 98] =  256;    assign rom_im[ 98] =    0;
      assign rom_re[ 99] =    0;    assign rom_im[ 99] = -256;
      assign rom_re[100] =  256;    assign rom_im[100] =    0;
      assign rom_re[101] =  181;    assign rom_im[101] = -181;
      assign rom_re[102] =  256;    assign rom_im[102] =    0;
      assign rom_re[103] = -181;    assign rom_im[103] = -181;
      assign rom_re[104] =  256;    assign rom_im[104] =    0;
      assign rom_re[105] =  256;    assign rom_im[105] =    0;
      assign rom_re[106] =  256;    assign rom_im[106] =    0;
      assign rom_re[107] =    0;    assign rom_im[107] = -256;
      assign rom_re[108] =  256;    assign rom_im[108] =    0;
      assign rom_re[109] =  181;    assign rom_im[109] = -181;
      assign rom_re[110] =  256;    assign rom_im[110] =    0;
      assign rom_re[111] = -181;    assign rom_im[111] = -181;
      assign rom_re[112] =  256;    assign rom_im[112] =    0;
      assign rom_re[113] =  256;    assign rom_im[113] =    0;
      assign rom_re[114] =  256;    assign rom_im[114] =    0;
      assign rom_re[115] =    0;    assign rom_im[115] = -256;
      assign rom_re[116] =  256;    assign rom_im[116] =    0;
      assign rom_re[117] =  181;    assign rom_im[117] = -181;
      assign rom_re[118] =  256;    assign rom_im[118] =    0;
      assign rom_re[119] = -181;    assign rom_im[119] = -181;
      assign rom_re[120] =  256;    assign rom_im[120] =    0;
      assign rom_re[121] =  256;    assign rom_im[121] =    0;
      assign rom_re[122] =  256;    assign rom_im[122] =    0;
      assign rom_re[123] =    0;    assign rom_im[123] = -256;
      assign rom_re[124] =  256;    assign rom_im[124] =    0;
      assign rom_re[125] =  181;    assign rom_im[125] = -181;
      assign rom_re[126] =  256;    assign rom_im[126] =    0;
      assign rom_re[127] = -181;    assign rom_im[127] = -181;
      assign rom_re[128] =  256;    assign rom_im[128] =    0;
      assign rom_re[129] =  256;    assign rom_im[129] =    0;
      assign rom_re[130] =  256;    assign rom_im[130] =    0;
      assign rom_re[131] =    0;    assign rom_im[131] = -256;
      assign rom_re[132] =  256;    assign rom_im[132] =    0;
      assign rom_re[133] =  181;    assign rom_im[133] = -181;
      assign rom_re[134] =  256;    assign rom_im[134] =    0;
      assign rom_re[135] = -181;    assign rom_im[135] = -181;
      assign rom_re[136] =  256;    assign rom_im[136] =    0;
      assign rom_re[137] =  256;    assign rom_im[137] =    0;
      assign rom_re[138] =  256;    assign rom_im[138] =    0;
      assign rom_re[139] =    0;    assign rom_im[139] = -256;
      assign rom_re[140] =  256;    assign rom_im[140] =    0;
      assign rom_re[141] =  181;    assign rom_im[141] = -181;
      assign rom_re[142] =  256;    assign rom_im[142] =    0;
      assign rom_re[143] = -181;    assign rom_im[143] = -181;
      assign rom_re[144] =  256;    assign rom_im[144] =    0;
      assign rom_re[145] =  256;    assign rom_im[145] =    0;
      assign rom_re[146] =  256;    assign rom_im[146] =    0;
      assign rom_re[147] =    0;    assign rom_im[147] = -256;
      assign rom_re[148] =  256;    assign rom_im[148] =    0;
      assign rom_re[149] =  181;    assign rom_im[149] = -181;
      assign rom_re[150] =  256;    assign rom_im[150] =    0;
      assign rom_re[151] = -181;    assign rom_im[151] = -181;
      assign rom_re[152] =  256;    assign rom_im[152] =    0;
      assign rom_re[153] =  256;    assign rom_im[153] =    0;
      assign rom_re[154] =  256;    assign rom_im[154] =    0;
      assign rom_re[155] =    0;    assign rom_im[155] = -256;
      assign rom_re[156] =  256;    assign rom_im[156] =    0;
      assign rom_re[157] =  181;    assign rom_im[157] = -181;
      assign rom_re[158] =  256;    assign rom_im[158] =    0;
      assign rom_re[159] = -181;    assign rom_im[159] = -181;
      assign rom_re[160] =  256;    assign rom_im[160] =    0;
      assign rom_re[161] =  256;    assign rom_im[161] =    0;
      assign rom_re[162] =  256;    assign rom_im[162] =    0;
      assign rom_re[163] =    0;    assign rom_im[163] = -256;
      assign rom_re[164] =  256;    assign rom_im[164] =    0;
      assign rom_re[165] =  181;    assign rom_im[165] = -181;
      assign rom_re[166] =  256;    assign rom_im[166] =    0;
      assign rom_re[167] = -181;    assign rom_im[167] = -181;
      assign rom_re[168] =  256;    assign rom_im[168] =    0;
      assign rom_re[169] =  256;    assign rom_im[169] =    0;
      assign rom_re[170] =  256;    assign rom_im[170] =    0;
      assign rom_re[171] =    0;    assign rom_im[171] = -256;
      assign rom_re[172] =  256;    assign rom_im[172] =    0;
      assign rom_re[173] =  181;    assign rom_im[173] = -181;
      assign rom_re[174] =  256;    assign rom_im[174] =    0;
      assign rom_re[175] = -181;    assign rom_im[175] = -181;
      assign rom_re[176] =  256;    assign rom_im[176] =    0;
      assign rom_re[177] =  256;    assign rom_im[177] =    0;
      assign rom_re[178] =  256;    assign rom_im[178] =    0;
      assign rom_re[179] =    0;    assign rom_im[179] = -256;
      assign rom_re[180] =  256;    assign rom_im[180] =    0;
      assign rom_re[181] =  181;    assign rom_im[181] = -181;
      assign rom_re[182] =  256;    assign rom_im[182] =    0;
      assign rom_re[183] = -181;    assign rom_im[183] = -181;
      assign rom_re[184] =  256;    assign rom_im[184] =    0;
      assign rom_re[185] =  256;    assign rom_im[185] =    0;
      assign rom_re[186] =  256;    assign rom_im[186] =    0;
      assign rom_re[187] =    0;    assign rom_im[187] = -256;
      assign rom_re[188] =  256;    assign rom_im[188] =    0;
      assign rom_re[189] =  181;    assign rom_im[189] = -181;
      assign rom_re[190] =  256;    assign rom_im[190] =    0;
      assign rom_re[191] = -181;    assign rom_im[191] = -181;
      assign rom_re[192] =  256;    assign rom_im[192] =    0;
      assign rom_re[193] =  256;    assign rom_im[193] =    0;
      assign rom_re[194] =  256;    assign rom_im[194] =    0;
      assign rom_re[195] =    0;    assign rom_im[195] = -256;
      assign rom_re[196] =  256;    assign rom_im[196] =    0;
      assign rom_re[197] =  181;    assign rom_im[197] = -181;
      assign rom_re[198] =  256;    assign rom_im[198] =    0;
      assign rom_re[199] = -181;    assign rom_im[199] = -181;
      assign rom_re[200] =  256;    assign rom_im[200] =    0;
      assign rom_re[201] =  256;    assign rom_im[201] =    0;
      assign rom_re[202] =  256;    assign rom_im[202] =    0;
      assign rom_re[203] =    0;    assign rom_im[203] = -256;
      assign rom_re[204] =  256;    assign rom_im[204] =    0;
      assign rom_re[205] =  181;    assign rom_im[205] = -181;
      assign rom_re[206] =  256;    assign rom_im[206] =    0;
      assign rom_re[207] = -181;    assign rom_im[207] = -181;
      assign rom_re[208] =  256;    assign rom_im[208] =    0;
      assign rom_re[209] =  256;    assign rom_im[209] =    0;
      assign rom_re[210] =  256;    assign rom_im[210] =    0;
      assign rom_re[211] =    0;    assign rom_im[211] = -256;
      assign rom_re[212] =  256;    assign rom_im[212] =    0;
      assign rom_re[213] =  181;    assign rom_im[213] = -181;
      assign rom_re[214] =  256;    assign rom_im[214] =    0;
      assign rom_re[215] = -181;    assign rom_im[215] = -181;
      assign rom_re[216] =  256;    assign rom_im[216] =    0;
      assign rom_re[217] =  256;    assign rom_im[217] =    0;
      assign rom_re[218] =  256;    assign rom_im[218] =    0;
      assign rom_re[219] =    0;    assign rom_im[219] = -256;
      assign rom_re[220] =  256;    assign rom_im[220] =    0;
      assign rom_re[221] =  181;    assign rom_im[221] = -181;
      assign rom_re[222] =  256;    assign rom_im[222] =    0;
      assign rom_re[223] = -181;    assign rom_im[223] = -181;
      assign rom_re[224] =  256;    assign rom_im[224] =    0;
      assign rom_re[225] =  256;    assign rom_im[225] =    0;
      assign rom_re[226] =  256;    assign rom_im[226] =    0;
      assign rom_re[227] =    0;    assign rom_im[227] = -256;
      assign rom_re[228] =  256;    assign rom_im[228] =    0;
      assign rom_re[229] =  181;    assign rom_im[229] = -181;
      assign rom_re[230] =  256;    assign rom_im[230] =    0;
      assign rom_re[231] = -181;    assign rom_im[231] = -181;
      assign rom_re[232] =  256;    assign rom_im[232] =    0;
      assign rom_re[233] =  256;    assign rom_im[233] =    0;
      assign rom_re[234] =  256;    assign rom_im[234] =    0;
      assign rom_re[235] =    0;    assign rom_im[235] = -256;
      assign rom_re[236] =  256;    assign rom_im[236] =    0;
      assign rom_re[237] =  181;    assign rom_im[237] = -181;
      assign rom_re[238] =  256;    assign rom_im[238] =    0;
      assign rom_re[239] = -181;    assign rom_im[239] = -181;
      assign rom_re[240] =  256;    assign rom_im[240] =    0;
      assign rom_re[241] =  256;    assign rom_im[241] =    0;
      assign rom_re[242] =  256;    assign rom_im[242] =    0;
      assign rom_re[243] =    0;    assign rom_im[243] = -256;
      assign rom_re[244] =  256;    assign rom_im[244] =    0;
      assign rom_re[245] =  181;    assign rom_im[245] = -181;
      assign rom_re[246] =  256;    assign rom_im[246] =    0;
      assign rom_re[247] = -181;    assign rom_im[247] = -181;
      assign rom_re[248] =  256;    assign rom_im[248] =    0;
      assign rom_re[249] =  256;    assign rom_im[249] =    0;
      assign rom_re[250] =  256;    assign rom_im[250] =    0;
      assign rom_re[251] =    0;    assign rom_im[251] = -256;
      assign rom_re[252] =  256;    assign rom_im[252] =    0;
      assign rom_re[253] =  181;    assign rom_im[253] = -181;
      assign rom_re[254] =  256;    assign rom_im[254] =    0;
      assign rom_re[255] = -181;    assign rom_im[255] = -181;
      assign rom_re[256] =  256;    assign rom_im[256] =    0;
      assign rom_re[257] =  256;    assign rom_im[257] =    0;
      assign rom_re[258] =  256;    assign rom_im[258] =    0;
      assign rom_re[259] =    0;    assign rom_im[259] = -256;
      assign rom_re[260] =  256;    assign rom_im[260] =    0;
      assign rom_re[261] =  181;    assign rom_im[261] = -181;
      assign rom_re[262] =  256;    assign rom_im[262] =    0;
      assign rom_re[263] = -181;    assign rom_im[263] = -181;
      assign rom_re[264] =  256;    assign rom_im[264] =    0;
      assign rom_re[265] =  256;    assign rom_im[265] =    0;
      assign rom_re[266] =  256;    assign rom_im[266] =    0;
      assign rom_re[267] =    0;    assign rom_im[267] = -256;
      assign rom_re[268] =  256;    assign rom_im[268] =    0;
      assign rom_re[269] =  181;    assign rom_im[269] = -181;
      assign rom_re[270] =  256;    assign rom_im[270] =    0;
      assign rom_re[271] = -181;    assign rom_im[271] = -181;
      assign rom_re[272] =  256;    assign rom_im[272] =    0;
      assign rom_re[273] =  256;    assign rom_im[273] =    0;
      assign rom_re[274] =  256;    assign rom_im[274] =    0;
      assign rom_re[275] =    0;    assign rom_im[275] = -256;
      assign rom_re[276] =  256;    assign rom_im[276] =    0;
      assign rom_re[277] =  181;    assign rom_im[277] = -181;
      assign rom_re[278] =  256;    assign rom_im[278] =    0;
      assign rom_re[279] = -181;    assign rom_im[279] = -181;
      assign rom_re[280] =  256;    assign rom_im[280] =    0;
      assign rom_re[281] =  256;    assign rom_im[281] =    0;
      assign rom_re[282] =  256;    assign rom_im[282] =    0;
      assign rom_re[283] =    0;    assign rom_im[283] = -256;
      assign rom_re[284] =  256;    assign rom_im[284] =    0;
      assign rom_re[285] =  181;    assign rom_im[285] = -181;
      assign rom_re[286] =  256;    assign rom_im[286] =    0;
      assign rom_re[287] = -181;    assign rom_im[287] = -181;
      assign rom_re[288] =  256;    assign rom_im[288] =    0;
      assign rom_re[289] =  256;    assign rom_im[289] =    0;
      assign rom_re[290] =  256;    assign rom_im[290] =    0;
      assign rom_re[291] =    0;    assign rom_im[291] = -256;
      assign rom_re[292] =  256;    assign rom_im[292] =    0;
      assign rom_re[293] =  181;    assign rom_im[293] = -181;
      assign rom_re[294] =  256;    assign rom_im[294] =    0;
      assign rom_re[295] = -181;    assign rom_im[295] = -181;
      assign rom_re[296] =  256;    assign rom_im[296] =    0;
      assign rom_re[297] =  256;    assign rom_im[297] =    0;
      assign rom_re[298] =  256;    assign rom_im[298] =    0;
      assign rom_re[299] =    0;    assign rom_im[299] = -256;
      assign rom_re[300] =  256;    assign rom_im[300] =    0;
      assign rom_re[301] =  181;    assign rom_im[301] = -181;
      assign rom_re[302] =  256;    assign rom_im[302] =    0;
      assign rom_re[303] = -181;    assign rom_im[303] = -181;
      assign rom_re[304] =  256;    assign rom_im[304] =    0;
      assign rom_re[305] =  256;    assign rom_im[305] =    0;
      assign rom_re[306] =  256;    assign rom_im[306] =    0;
      assign rom_re[307] =    0;    assign rom_im[307] = -256;
      assign rom_re[308] =  256;    assign rom_im[308] =    0;
      assign rom_re[309] =  181;    assign rom_im[309] = -181;
      assign rom_re[310] =  256;    assign rom_im[310] =    0;
      assign rom_re[311] = -181;    assign rom_im[311] = -181;
      assign rom_re[312] =  256;    assign rom_im[312] =    0;
      assign rom_re[313] =  256;    assign rom_im[313] =    0;
      assign rom_re[314] =  256;    assign rom_im[314] =    0;
      assign rom_re[315] =    0;    assign rom_im[315] = -256;
      assign rom_re[316] =  256;    assign rom_im[316] =    0;
      assign rom_re[317] =  181;    assign rom_im[317] = -181;
      assign rom_re[318] =  256;    assign rom_im[318] =    0;
      assign rom_re[319] = -181;    assign rom_im[319] = -181;
      assign rom_re[320] =  256;    assign rom_im[320] =    0;
      assign rom_re[321] =  256;    assign rom_im[321] =    0;
      assign rom_re[322] =  256;    assign rom_im[322] =    0;
      assign rom_re[323] =    0;    assign rom_im[323] = -256;
      assign rom_re[324] =  256;    assign rom_im[324] =    0;
      assign rom_re[325] =  181;    assign rom_im[325] = -181;
      assign rom_re[326] =  256;    assign rom_im[326] =    0;
      assign rom_re[327] = -181;    assign rom_im[327] = -181;
      assign rom_re[328] =  256;    assign rom_im[328] =    0;
      assign rom_re[329] =  256;    assign rom_im[329] =    0;
      assign rom_re[330] =  256;    assign rom_im[330] =    0;
      assign rom_re[331] =    0;    assign rom_im[331] = -256;
      assign rom_re[332] =  256;    assign rom_im[332] =    0;
      assign rom_re[333] =  181;    assign rom_im[333] = -181;
      assign rom_re[334] =  256;    assign rom_im[334] =    0;
      assign rom_re[335] = -181;    assign rom_im[335] = -181;
      assign rom_re[336] =  256;    assign rom_im[336] =    0;
      assign rom_re[337] =  256;    assign rom_im[337] =    0;
      assign rom_re[338] =  256;    assign rom_im[338] =    0;
      assign rom_re[339] =    0;    assign rom_im[339] = -256;
      assign rom_re[340] =  256;    assign rom_im[340] =    0;
      assign rom_re[341] =  181;    assign rom_im[341] = -181;
      assign rom_re[342] =  256;    assign rom_im[342] =    0;
      assign rom_re[343] = -181;    assign rom_im[343] = -181;
      assign rom_re[344] =  256;    assign rom_im[344] =    0;
      assign rom_re[345] =  256;    assign rom_im[345] =    0;
      assign rom_re[346] =  256;    assign rom_im[346] =    0;
      assign rom_re[347] =    0;    assign rom_im[347] = -256;
      assign rom_re[348] =  256;    assign rom_im[348] =    0;
      assign rom_re[349] =  181;    assign rom_im[349] = -181;
      assign rom_re[350] =  256;    assign rom_im[350] =    0;
      assign rom_re[351] = -181;    assign rom_im[351] = -181;
      assign rom_re[352] =  256;    assign rom_im[352] =    0;
      assign rom_re[353] =  256;    assign rom_im[353] =    0;
      assign rom_re[354] =  256;    assign rom_im[354] =    0;
      assign rom_re[355] =    0;    assign rom_im[355] = -256;
      assign rom_re[356] =  256;    assign rom_im[356] =    0;
      assign rom_re[357] =  181;    assign rom_im[357] = -181;
      assign rom_re[358] =  256;    assign rom_im[358] =    0;
      assign rom_re[359] = -181;    assign rom_im[359] = -181;
      assign rom_re[360] =  256;    assign rom_im[360] =    0;
      assign rom_re[361] =  256;    assign rom_im[361] =    0;
      assign rom_re[362] =  256;    assign rom_im[362] =    0;
      assign rom_re[363] =    0;    assign rom_im[363] = -256;
      assign rom_re[364] =  256;    assign rom_im[364] =    0;
      assign rom_re[365] =  181;    assign rom_im[365] = -181;
      assign rom_re[366] =  256;    assign rom_im[366] =    0;
      assign rom_re[367] = -181;    assign rom_im[367] = -181;
      assign rom_re[368] =  256;    assign rom_im[368] =    0;
      assign rom_re[369] =  256;    assign rom_im[369] =    0;
      assign rom_re[370] =  256;    assign rom_im[370] =    0;
      assign rom_re[371] =    0;    assign rom_im[371] = -256;
      assign rom_re[372] =  256;    assign rom_im[372] =    0;
      assign rom_re[373] =  181;    assign rom_im[373] = -181;
      assign rom_re[374] =  256;    assign rom_im[374] =    0;
      assign rom_re[375] = -181;    assign rom_im[375] = -181;
      assign rom_re[376] =  256;    assign rom_im[376] =    0;
      assign rom_re[377] =  256;    assign rom_im[377] =    0;
      assign rom_re[378] =  256;    assign rom_im[378] =    0;
      assign rom_re[379] =    0;    assign rom_im[379] = -256;
      assign rom_re[380] =  256;    assign rom_im[380] =    0;
      assign rom_re[381] =  181;    assign rom_im[381] = -181;
      assign rom_re[382] =  256;    assign rom_im[382] =    0;
      assign rom_re[383] = -181;    assign rom_im[383] = -181;
      assign rom_re[384] =  256;    assign rom_im[384] =    0;
      assign rom_re[385] =  256;    assign rom_im[385] =    0;
      assign rom_re[386] =  256;    assign rom_im[386] =    0;
      assign rom_re[387] =    0;    assign rom_im[387] = -256;
      assign rom_re[388] =  256;    assign rom_im[388] =    0;
      assign rom_re[389] =  181;    assign rom_im[389] = -181;
      assign rom_re[390] =  256;    assign rom_im[390] =    0;
      assign rom_re[391] = -181;    assign rom_im[391] = -181;
      assign rom_re[392] =  256;    assign rom_im[392] =    0;
      assign rom_re[393] =  256;    assign rom_im[393] =    0;
      assign rom_re[394] =  256;    assign rom_im[394] =    0;
      assign rom_re[395] =    0;    assign rom_im[395] = -256;
      assign rom_re[396] =  256;    assign rom_im[396] =    0;
      assign rom_re[397] =  181;    assign rom_im[397] = -181;
      assign rom_re[398] =  256;    assign rom_im[398] =    0;
      assign rom_re[399] = -181;    assign rom_im[399] = -181;
      assign rom_re[400] =  256;    assign rom_im[400] =    0;
      assign rom_re[401] =  256;    assign rom_im[401] =    0;
      assign rom_re[402] =  256;    assign rom_im[402] =    0;
      assign rom_re[403] =    0;    assign rom_im[403] = -256;
      assign rom_re[404] =  256;    assign rom_im[404] =    0;
      assign rom_re[405] =  181;    assign rom_im[405] = -181;
      assign rom_re[406] =  256;    assign rom_im[406] =    0;
      assign rom_re[407] = -181;    assign rom_im[407] = -181;
      assign rom_re[408] =  256;    assign rom_im[408] =    0;
      assign rom_re[409] =  256;    assign rom_im[409] =    0;
      assign rom_re[410] =  256;    assign rom_im[410] =    0;
      assign rom_re[411] =    0;    assign rom_im[411] = -256;
      assign rom_re[412] =  256;    assign rom_im[412] =    0;
      assign rom_re[413] =  181;    assign rom_im[413] = -181;
      assign rom_re[414] =  256;    assign rom_im[414] =    0;
      assign rom_re[415] = -181;    assign rom_im[415] = -181;
      assign rom_re[416] =  256;    assign rom_im[416] =    0;
      assign rom_re[417] =  256;    assign rom_im[417] =    0;
      assign rom_re[418] =  256;    assign rom_im[418] =    0;
      assign rom_re[419] =    0;    assign rom_im[419] = -256;
      assign rom_re[420] =  256;    assign rom_im[420] =    0;
      assign rom_re[421] =  181;    assign rom_im[421] = -181;
      assign rom_re[422] =  256;    assign rom_im[422] =    0;
      assign rom_re[423] = -181;    assign rom_im[423] = -181;
      assign rom_re[424] =  256;    assign rom_im[424] =    0;
      assign rom_re[425] =  256;    assign rom_im[425] =    0;
      assign rom_re[426] =  256;    assign rom_im[426] =    0;
      assign rom_re[427] =    0;    assign rom_im[427] = -256;
      assign rom_re[428] =  256;    assign rom_im[428] =    0;
      assign rom_re[429] =  181;    assign rom_im[429] = -181;
      assign rom_re[430] =  256;    assign rom_im[430] =    0;
      assign rom_re[431] = -181;    assign rom_im[431] = -181;
      assign rom_re[432] =  256;    assign rom_im[432] =    0;
      assign rom_re[433] =  256;    assign rom_im[433] =    0;
      assign rom_re[434] =  256;    assign rom_im[434] =    0;
      assign rom_re[435] =    0;    assign rom_im[435] = -256;
      assign rom_re[436] =  256;    assign rom_im[436] =    0;
      assign rom_re[437] =  181;    assign rom_im[437] = -181;
      assign rom_re[438] =  256;    assign rom_im[438] =    0;
      assign rom_re[439] = -181;    assign rom_im[439] = -181;
      assign rom_re[440] =  256;    assign rom_im[440] =    0;
      assign rom_re[441] =  256;    assign rom_im[441] =    0;
      assign rom_re[442] =  256;    assign rom_im[442] =    0;
      assign rom_re[443] =    0;    assign rom_im[443] = -256;
      assign rom_re[444] =  256;    assign rom_im[444] =    0;
      assign rom_re[445] =  181;    assign rom_im[445] = -181;
      assign rom_re[446] =  256;    assign rom_im[446] =    0;
      assign rom_re[447] = -181;    assign rom_im[447] = -181;
      assign rom_re[448] =  256;    assign rom_im[448] =    0;
      assign rom_re[449] =  256;    assign rom_im[449] =    0;
      assign rom_re[450] =  256;    assign rom_im[450] =    0;
      assign rom_re[451] =    0;    assign rom_im[451] = -256;
      assign rom_re[452] =  256;    assign rom_im[452] =    0;
      assign rom_re[453] =  181;    assign rom_im[453] = -181;
      assign rom_re[454] =  256;    assign rom_im[454] =    0;
      assign rom_re[455] = -181;    assign rom_im[455] = -181;
      assign rom_re[456] =  256;    assign rom_im[456] =    0;
      assign rom_re[457] =  256;    assign rom_im[457] =    0;
      assign rom_re[458] =  256;    assign rom_im[458] =    0;
      assign rom_re[459] =    0;    assign rom_im[459] = -256;
      assign rom_re[460] =  256;    assign rom_im[460] =    0;
      assign rom_re[461] =  181;    assign rom_im[461] = -181;
      assign rom_re[462] =  256;    assign rom_im[462] =    0;
      assign rom_re[463] = -181;    assign rom_im[463] = -181;
      assign rom_re[464] =  256;    assign rom_im[464] =    0;
      assign rom_re[465] =  256;    assign rom_im[465] =    0;
      assign rom_re[466] =  256;    assign rom_im[466] =    0;
      assign rom_re[467] =    0;    assign rom_im[467] = -256;
      assign rom_re[468] =  256;    assign rom_im[468] =    0;
      assign rom_re[469] =  181;    assign rom_im[469] = -181;
      assign rom_re[470] =  256;    assign rom_im[470] =    0;
      assign rom_re[471] = -181;    assign rom_im[471] = -181;
      assign rom_re[472] =  256;    assign rom_im[472] =    0;
      assign rom_re[473] =  256;    assign rom_im[473] =    0;
      assign rom_re[474] =  256;    assign rom_im[474] =    0;
      assign rom_re[475] =    0;    assign rom_im[475] = -256;
      assign rom_re[476] =  256;    assign rom_im[476] =    0;
      assign rom_re[477] =  181;    assign rom_im[477] = -181;
      assign rom_re[478] =  256;    assign rom_im[478] =    0;
      assign rom_re[479] = -181;    assign rom_im[479] = -181;
      assign rom_re[480] =  256;    assign rom_im[480] =    0;
      assign rom_re[481] =  256;    assign rom_im[481] =    0;
      assign rom_re[482] =  256;    assign rom_im[482] =    0;
      assign rom_re[483] =    0;    assign rom_im[483] = -256;
      assign rom_re[484] =  256;    assign rom_im[484] =    0;
      assign rom_re[485] =  181;    assign rom_im[485] = -181;
      assign rom_re[486] =  256;    assign rom_im[486] =    0;
      assign rom_re[487] = -181;    assign rom_im[487] = -181;
      assign rom_re[488] =  256;    assign rom_im[488] =    0;
      assign rom_re[489] =  256;    assign rom_im[489] =    0;
      assign rom_re[490] =  256;    assign rom_im[490] =    0;
      assign rom_re[491] =    0;    assign rom_im[491] = -256;
      assign rom_re[492] =  256;    assign rom_im[492] =    0;
      assign rom_re[493] =  181;    assign rom_im[493] = -181;
      assign rom_re[494] =  256;    assign rom_im[494] =    0;
      assign rom_re[495] = -181;    assign rom_im[495] = -181;
      assign rom_re[496] =  256;    assign rom_im[496] =    0;
      assign rom_re[497] =  256;    assign rom_im[497] =    0;
      assign rom_re[498] =  256;    assign rom_im[498] =    0;
      assign rom_re[499] =    0;    assign rom_im[499] = -256;
      assign rom_re[500] =  256;    assign rom_im[500] =    0;
      assign rom_re[501] =  181;    assign rom_im[501] = -181;
      assign rom_re[502] =  256;    assign rom_im[502] =    0;
      assign rom_re[503] = -181;    assign rom_im[503] = -181;
      assign rom_re[504] =  256;    assign rom_im[504] =    0;
      assign rom_re[505] =  256;    assign rom_im[505] =    0;
      assign rom_re[506] =  256;    assign rom_im[506] =    0;
      assign rom_re[507] =    0;    assign rom_im[507] = -256;
      assign rom_re[508] =  256;    assign rom_im[508] =    0;
      assign rom_re[509] =  181;    assign rom_im[509] = -181;
      assign rom_re[510] =  256;    assign rom_im[510] =    0;
      assign rom_re[511] = -181;    assign rom_im[511] = -181;

     endmodule
